module DRAM (
input wire [15:0] address,
input clock,
input wire [7:0] data,
input wren,
output reg [7:0] q);
reg [7:0] DRAM[131071:0];

initial begin
DRAM[0] = 8'b10100001;
DRAM[1] = 8'b10011111;
DRAM[2] = 8'b10100000;
DRAM[3] = 8'b10011111;
DRAM[4] = 8'b10011110;
DRAM[5] = 8'b10011100;
DRAM[6] = 8'b10011010;
DRAM[7] = 8'b10011011;
DRAM[8] = 8'b10011110;
DRAM[9] = 8'b10100110;
DRAM[10] = 8'b10101000;
DRAM[11] = 8'b10101100;
DRAM[12] = 8'b10101101;
DRAM[13] = 8'b10100100;
DRAM[14] = 8'b10010000;
DRAM[15] = 8'b01110000;
DRAM[16] = 8'b01011110;
DRAM[17] = 8'b01100000;
DRAM[18] = 8'b01100111;
DRAM[19] = 8'b01101011;
DRAM[20] = 8'b01101011;
DRAM[21] = 8'b01101101;
DRAM[22] = 8'b01101011;
DRAM[23] = 8'b01101101;
DRAM[24] = 8'b01101101;
DRAM[25] = 8'b01101011;
DRAM[26] = 8'b01101110;
DRAM[27] = 8'b01110110;
DRAM[28] = 8'b01111010;
DRAM[29] = 8'b01111011;
DRAM[30] = 8'b01111110;
DRAM[31] = 8'b10000001;
DRAM[32] = 8'b10000001;
DRAM[33] = 8'b10000000;
DRAM[34] = 8'b10000111;
DRAM[35] = 8'b10000010;
DRAM[36] = 8'b01111110;
DRAM[37] = 8'b10000010;
DRAM[38] = 8'b10000010;
DRAM[39] = 8'b10000110;
DRAM[40] = 8'b10000110;
DRAM[41] = 8'b10000110;
DRAM[42] = 8'b10001000;
DRAM[43] = 8'b10000100;
DRAM[44] = 8'b10000101;
DRAM[45] = 8'b10000100;
DRAM[46] = 8'b10000111;
DRAM[47] = 8'b10000011;
DRAM[48] = 8'b10000111;
DRAM[49] = 8'b10001010;
DRAM[50] = 8'b10000110;
DRAM[51] = 8'b10000110;
DRAM[52] = 8'b10000111;
DRAM[53] = 8'b10000011;
DRAM[54] = 8'b10000001;
DRAM[55] = 8'b10000011;
DRAM[56] = 8'b10000011;
DRAM[57] = 8'b10000110;
DRAM[58] = 8'b10000100;
DRAM[59] = 8'b10000100;
DRAM[60] = 8'b10000110;
DRAM[61] = 8'b10001000;
DRAM[62] = 8'b10000101;
DRAM[63] = 8'b10000101;
DRAM[64] = 8'b10001001;
DRAM[65] = 8'b10000001;
DRAM[66] = 8'b10000100;
DRAM[67] = 8'b10000011;
DRAM[68] = 8'b10000001;
DRAM[69] = 8'b10000100;
DRAM[70] = 8'b10000001;
DRAM[71] = 8'b10000001;
DRAM[72] = 8'b10000010;
DRAM[73] = 8'b01111110;
DRAM[74] = 8'b10000001;
DRAM[75] = 8'b10000010;
DRAM[76] = 8'b01111010;
DRAM[77] = 8'b01111000;
DRAM[78] = 8'b01110001;
DRAM[79] = 8'b01101000;
DRAM[80] = 8'b01110011;
DRAM[81] = 8'b10000111;
DRAM[82] = 8'b10010011;
DRAM[83] = 8'b10011011;
DRAM[84] = 8'b10011110;
DRAM[85] = 8'b10011110;
DRAM[86] = 8'b10010110;
DRAM[87] = 8'b10011001;
DRAM[88] = 8'b10011011;
DRAM[89] = 8'b10011010;
DRAM[90] = 8'b10011101;
DRAM[91] = 8'b10011011;
DRAM[92] = 8'b10010111;
DRAM[93] = 8'b10011001;
DRAM[94] = 8'b10011010;
DRAM[95] = 8'b10011001;
DRAM[96] = 8'b10011101;
DRAM[97] = 8'b10011011;
DRAM[98] = 8'b10011111;
DRAM[99] = 8'b10011010;
DRAM[100] = 8'b10100110;
DRAM[101] = 8'b11001011;
DRAM[102] = 8'b11010110;
DRAM[103] = 8'b11011010;
DRAM[104] = 8'b11010001;
DRAM[105] = 8'b10010010;
DRAM[106] = 8'b01101000;
DRAM[107] = 8'b01110000;
DRAM[108] = 8'b01110100;
DRAM[109] = 8'b01111000;
DRAM[110] = 8'b01110111;
DRAM[111] = 8'b01111001;
DRAM[112] = 8'b01111110;
DRAM[113] = 8'b01110110;
DRAM[114] = 8'b01111001;
DRAM[115] = 8'b01111010;
DRAM[116] = 8'b01111001;
DRAM[117] = 8'b01111110;
DRAM[118] = 8'b01111101;
DRAM[119] = 8'b01111001;
DRAM[120] = 8'b01111100;
DRAM[121] = 8'b10000000;
DRAM[122] = 8'b01111010;
DRAM[123] = 8'b01111100;
DRAM[124] = 8'b01111000;
DRAM[125] = 8'b01110111;
DRAM[126] = 8'b10101000;
DRAM[127] = 8'b10010100;
DRAM[128] = 8'b10011110;
DRAM[129] = 8'b10011110;
DRAM[130] = 8'b10011111;
DRAM[131] = 8'b10011001;
DRAM[132] = 8'b10011011;
DRAM[133] = 8'b10011000;
DRAM[134] = 8'b10011010;
DRAM[135] = 8'b10011001;
DRAM[136] = 8'b10011001;
DRAM[137] = 8'b10100000;
DRAM[138] = 8'b10101001;
DRAM[139] = 8'b10101100;
DRAM[140] = 8'b10101101;
DRAM[141] = 8'b10100000;
DRAM[142] = 8'b10001100;
DRAM[143] = 8'b01110011;
DRAM[144] = 8'b01011100;
DRAM[145] = 8'b01011100;
DRAM[146] = 8'b01100100;
DRAM[147] = 8'b01101011;
DRAM[148] = 8'b01101000;
DRAM[149] = 8'b01101010;
DRAM[150] = 8'b01100110;
DRAM[151] = 8'b01101001;
DRAM[152] = 8'b01101000;
DRAM[153] = 8'b01101000;
DRAM[154] = 8'b01101111;
DRAM[155] = 8'b01110101;
DRAM[156] = 8'b01111010;
DRAM[157] = 8'b01111110;
DRAM[158] = 8'b01111100;
DRAM[159] = 8'b01111100;
DRAM[160] = 8'b10000011;
DRAM[161] = 8'b10000000;
DRAM[162] = 8'b10000011;
DRAM[163] = 8'b10000010;
DRAM[164] = 8'b10000010;
DRAM[165] = 8'b10000100;
DRAM[166] = 8'b10000010;
DRAM[167] = 8'b10000101;
DRAM[168] = 8'b10000110;
DRAM[169] = 8'b10000111;
DRAM[170] = 8'b10000101;
DRAM[171] = 8'b10000101;
DRAM[172] = 8'b10000101;
DRAM[173] = 8'b10000100;
DRAM[174] = 8'b10000010;
DRAM[175] = 8'b10000100;
DRAM[176] = 8'b10000110;
DRAM[177] = 8'b10000100;
DRAM[178] = 8'b10000011;
DRAM[179] = 8'b10000100;
DRAM[180] = 8'b10000110;
DRAM[181] = 8'b10000010;
DRAM[182] = 8'b10000010;
DRAM[183] = 8'b10000010;
DRAM[184] = 8'b10000011;
DRAM[185] = 8'b10000010;
DRAM[186] = 8'b10000001;
DRAM[187] = 8'b10000011;
DRAM[188] = 8'b10000110;
DRAM[189] = 8'b10000010;
DRAM[190] = 8'b10000010;
DRAM[191] = 8'b10000100;
DRAM[192] = 8'b10000110;
DRAM[193] = 8'b10000001;
DRAM[194] = 8'b10000000;
DRAM[195] = 8'b10000010;
DRAM[196] = 8'b10000000;
DRAM[197] = 8'b10000010;
DRAM[198] = 8'b10000000;
DRAM[199] = 8'b10000000;
DRAM[200] = 8'b10000001;
DRAM[201] = 8'b10000010;
DRAM[202] = 8'b10000010;
DRAM[203] = 8'b01111100;
DRAM[204] = 8'b01111000;
DRAM[205] = 8'b01110111;
DRAM[206] = 8'b01110001;
DRAM[207] = 8'b01101010;
DRAM[208] = 8'b01110000;
DRAM[209] = 8'b10000011;
DRAM[210] = 8'b10010001;
DRAM[211] = 8'b10011001;
DRAM[212] = 8'b10100001;
DRAM[213] = 8'b10011100;
DRAM[214] = 8'b10011001;
DRAM[215] = 8'b10011000;
DRAM[216] = 8'b10011000;
DRAM[217] = 8'b10011001;
DRAM[218] = 8'b10011010;
DRAM[219] = 8'b10011001;
DRAM[220] = 8'b10011000;
DRAM[221] = 8'b10011000;
DRAM[222] = 8'b10011011;
DRAM[223] = 8'b10011001;
DRAM[224] = 8'b10011001;
DRAM[225] = 8'b10011011;
DRAM[226] = 8'b10011100;
DRAM[227] = 8'b10011001;
DRAM[228] = 8'b10011011;
DRAM[229] = 8'b11000100;
DRAM[230] = 8'b11010100;
DRAM[231] = 8'b11011001;
DRAM[232] = 8'b11010111;
DRAM[233] = 8'b10110000;
DRAM[234] = 8'b01101010;
DRAM[235] = 8'b01101010;
DRAM[236] = 8'b01110100;
DRAM[237] = 8'b01110110;
DRAM[238] = 8'b01111000;
DRAM[239] = 8'b01111000;
DRAM[240] = 8'b01111010;
DRAM[241] = 8'b01111010;
DRAM[242] = 8'b01111010;
DRAM[243] = 8'b01111100;
DRAM[244] = 8'b01111100;
DRAM[245] = 8'b01111100;
DRAM[246] = 8'b01111101;
DRAM[247] = 8'b01111000;
DRAM[248] = 8'b01111011;
DRAM[249] = 8'b01111111;
DRAM[250] = 8'b01111110;
DRAM[251] = 8'b01111101;
DRAM[252] = 8'b01111010;
DRAM[253] = 8'b01111100;
DRAM[254] = 8'b01101111;
DRAM[255] = 8'b01000101;
DRAM[256] = 8'b10011101;
DRAM[257] = 8'b10011001;
DRAM[258] = 8'b10011100;
DRAM[259] = 8'b10011011;
DRAM[260] = 8'b10011011;
DRAM[261] = 8'b10011011;
DRAM[262] = 8'b10011001;
DRAM[263] = 8'b10011010;
DRAM[264] = 8'b10011101;
DRAM[265] = 8'b10100100;
DRAM[266] = 8'b10101001;
DRAM[267] = 8'b10101100;
DRAM[268] = 8'b10101001;
DRAM[269] = 8'b10011101;
DRAM[270] = 8'b10000111;
DRAM[271] = 8'b01110000;
DRAM[272] = 8'b01011100;
DRAM[273] = 8'b01011010;
DRAM[274] = 8'b01100001;
DRAM[275] = 8'b01100101;
DRAM[276] = 8'b01100110;
DRAM[277] = 8'b01101011;
DRAM[278] = 8'b01101000;
DRAM[279] = 8'b01100111;
DRAM[280] = 8'b01101000;
DRAM[281] = 8'b01101011;
DRAM[282] = 8'b01101111;
DRAM[283] = 8'b01110011;
DRAM[284] = 8'b01110110;
DRAM[285] = 8'b01111010;
DRAM[286] = 8'b01111101;
DRAM[287] = 8'b01111110;
DRAM[288] = 8'b10000000;
DRAM[289] = 8'b10000000;
DRAM[290] = 8'b10000000;
DRAM[291] = 8'b10000001;
DRAM[292] = 8'b10000010;
DRAM[293] = 8'b10000010;
DRAM[294] = 8'b10000011;
DRAM[295] = 8'b10000011;
DRAM[296] = 8'b10000010;
DRAM[297] = 8'b10000101;
DRAM[298] = 8'b10000101;
DRAM[299] = 8'b10000101;
DRAM[300] = 8'b10000011;
DRAM[301] = 8'b10000100;
DRAM[302] = 8'b10000110;
DRAM[303] = 8'b10000110;
DRAM[304] = 8'b10000011;
DRAM[305] = 8'b10000001;
DRAM[306] = 8'b10000011;
DRAM[307] = 8'b10000010;
DRAM[308] = 8'b10000011;
DRAM[309] = 8'b10000001;
DRAM[310] = 8'b10000000;
DRAM[311] = 8'b10000001;
DRAM[312] = 8'b10000010;
DRAM[313] = 8'b10000010;
DRAM[314] = 8'b10000001;
DRAM[315] = 8'b10000010;
DRAM[316] = 8'b10000100;
DRAM[317] = 8'b10000100;
DRAM[318] = 8'b10000100;
DRAM[319] = 8'b10000000;
DRAM[320] = 8'b10000010;
DRAM[321] = 8'b10000010;
DRAM[322] = 8'b10000001;
DRAM[323] = 8'b01111111;
DRAM[324] = 8'b01111111;
DRAM[325] = 8'b10000000;
DRAM[326] = 8'b10000000;
DRAM[327] = 8'b10000000;
DRAM[328] = 8'b01111110;
DRAM[329] = 8'b01111111;
DRAM[330] = 8'b01111111;
DRAM[331] = 8'b01111111;
DRAM[332] = 8'b01111100;
DRAM[333] = 8'b01111000;
DRAM[334] = 8'b01110010;
DRAM[335] = 8'b01101110;
DRAM[336] = 8'b01101011;
DRAM[337] = 8'b01110100;
DRAM[338] = 8'b10001000;
DRAM[339] = 8'b10010011;
DRAM[340] = 8'b10011100;
DRAM[341] = 8'b10011110;
DRAM[342] = 8'b10011010;
DRAM[343] = 8'b10011011;
DRAM[344] = 8'b10011110;
DRAM[345] = 8'b10011101;
DRAM[346] = 8'b10011010;
DRAM[347] = 8'b10011100;
DRAM[348] = 8'b10011011;
DRAM[349] = 8'b10011000;
DRAM[350] = 8'b10011010;
DRAM[351] = 8'b10011000;
DRAM[352] = 8'b10011010;
DRAM[353] = 8'b10011010;
DRAM[354] = 8'b10011011;
DRAM[355] = 8'b10010110;
DRAM[356] = 8'b10011000;
DRAM[357] = 8'b10101000;
DRAM[358] = 8'b11001101;
DRAM[359] = 8'b11010111;
DRAM[360] = 8'b11011010;
DRAM[361] = 8'b11001101;
DRAM[362] = 8'b10001100;
DRAM[363] = 8'b01101001;
DRAM[364] = 8'b01101111;
DRAM[365] = 8'b01110100;
DRAM[366] = 8'b01111001;
DRAM[367] = 8'b01110111;
DRAM[368] = 8'b01111011;
DRAM[369] = 8'b01111001;
DRAM[370] = 8'b01111000;
DRAM[371] = 8'b01111010;
DRAM[372] = 8'b01111010;
DRAM[373] = 8'b01111010;
DRAM[374] = 8'b01111101;
DRAM[375] = 8'b01111100;
DRAM[376] = 8'b01111101;
DRAM[377] = 8'b01111101;
DRAM[378] = 8'b01111110;
DRAM[379] = 8'b10000001;
DRAM[380] = 8'b10000000;
DRAM[381] = 8'b01011010;
DRAM[382] = 8'b00101111;
DRAM[383] = 8'b00101110;
DRAM[384] = 8'b10011101;
DRAM[385] = 8'b10011100;
DRAM[386] = 8'b10011101;
DRAM[387] = 8'b10011100;
DRAM[388] = 8'b10011011;
DRAM[389] = 8'b10011100;
DRAM[390] = 8'b10011100;
DRAM[391] = 8'b10011101;
DRAM[392] = 8'b10100011;
DRAM[393] = 8'b10100111;
DRAM[394] = 8'b10101001;
DRAM[395] = 8'b10101001;
DRAM[396] = 8'b10100011;
DRAM[397] = 8'b10011001;
DRAM[398] = 8'b10001000;
DRAM[399] = 8'b01110000;
DRAM[400] = 8'b01011010;
DRAM[401] = 8'b01011010;
DRAM[402] = 8'b01100100;
DRAM[403] = 8'b01100110;
DRAM[404] = 8'b01101010;
DRAM[405] = 8'b01101010;
DRAM[406] = 8'b01101001;
DRAM[407] = 8'b01100111;
DRAM[408] = 8'b01100111;
DRAM[409] = 8'b01101010;
DRAM[410] = 8'b01101111;
DRAM[411] = 8'b01110011;
DRAM[412] = 8'b01110110;
DRAM[413] = 8'b01111010;
DRAM[414] = 8'b01111100;
DRAM[415] = 8'b01111110;
DRAM[416] = 8'b10000000;
DRAM[417] = 8'b10000001;
DRAM[418] = 8'b10000001;
DRAM[419] = 8'b10000011;
DRAM[420] = 8'b10000011;
DRAM[421] = 8'b10000011;
DRAM[422] = 8'b10000001;
DRAM[423] = 8'b10000011;
DRAM[424] = 8'b10000101;
DRAM[425] = 8'b10000101;
DRAM[426] = 8'b10000100;
DRAM[427] = 8'b10000110;
DRAM[428] = 8'b10000100;
DRAM[429] = 8'b10000101;
DRAM[430] = 8'b10000101;
DRAM[431] = 8'b10000100;
DRAM[432] = 8'b10000101;
DRAM[433] = 8'b10000010;
DRAM[434] = 8'b10000010;
DRAM[435] = 8'b10000010;
DRAM[436] = 8'b10000100;
DRAM[437] = 8'b10000011;
DRAM[438] = 8'b10000010;
DRAM[439] = 8'b10000001;
DRAM[440] = 8'b10000010;
DRAM[441] = 8'b10000011;
DRAM[442] = 8'b10000000;
DRAM[443] = 8'b10000100;
DRAM[444] = 8'b10000101;
DRAM[445] = 8'b10000110;
DRAM[446] = 8'b10000010;
DRAM[447] = 8'b10000100;
DRAM[448] = 8'b10000011;
DRAM[449] = 8'b10000010;
DRAM[450] = 8'b10000110;
DRAM[451] = 8'b10000001;
DRAM[452] = 8'b10000000;
DRAM[453] = 8'b10000000;
DRAM[454] = 8'b10000000;
DRAM[455] = 8'b10000011;
DRAM[456] = 8'b01111110;
DRAM[457] = 8'b10000001;
DRAM[458] = 8'b10000010;
DRAM[459] = 8'b10000001;
DRAM[460] = 8'b01111110;
DRAM[461] = 8'b01111001;
DRAM[462] = 8'b01110001;
DRAM[463] = 8'b01101111;
DRAM[464] = 8'b01101100;
DRAM[465] = 8'b01101101;
DRAM[466] = 8'b10000100;
DRAM[467] = 8'b10010010;
DRAM[468] = 8'b10011001;
DRAM[469] = 8'b10011111;
DRAM[470] = 8'b10100000;
DRAM[471] = 8'b10011110;
DRAM[472] = 8'b10011110;
DRAM[473] = 8'b10100001;
DRAM[474] = 8'b10100001;
DRAM[475] = 8'b10011110;
DRAM[476] = 8'b10011101;
DRAM[477] = 8'b10011011;
DRAM[478] = 8'b10011010;
DRAM[479] = 8'b10011011;
DRAM[480] = 8'b10011010;
DRAM[481] = 8'b10011000;
DRAM[482] = 8'b10011000;
DRAM[483] = 8'b10010111;
DRAM[484] = 8'b10010111;
DRAM[485] = 8'b10010110;
DRAM[486] = 8'b10111101;
DRAM[487] = 8'b11010011;
DRAM[488] = 8'b11011010;
DRAM[489] = 8'b11011011;
DRAM[490] = 8'b10111011;
DRAM[491] = 8'b01110011;
DRAM[492] = 8'b01101111;
DRAM[493] = 8'b01110000;
DRAM[494] = 8'b01110111;
DRAM[495] = 8'b01110111;
DRAM[496] = 8'b01111000;
DRAM[497] = 8'b01111011;
DRAM[498] = 8'b01111000;
DRAM[499] = 8'b01111011;
DRAM[500] = 8'b01111000;
DRAM[501] = 8'b01111010;
DRAM[502] = 8'b01111100;
DRAM[503] = 8'b01111010;
DRAM[504] = 8'b01111111;
DRAM[505] = 8'b10000000;
DRAM[506] = 8'b10000011;
DRAM[507] = 8'b10000001;
DRAM[508] = 8'b01011000;
DRAM[509] = 8'b00110101;
DRAM[510] = 8'b00101100;
DRAM[511] = 8'b00110001;
DRAM[512] = 8'b10011100;
DRAM[513] = 8'b10011011;
DRAM[514] = 8'b10011101;
DRAM[515] = 8'b10011100;
DRAM[516] = 8'b10011100;
DRAM[517] = 8'b10011100;
DRAM[518] = 8'b10011000;
DRAM[519] = 8'b10011111;
DRAM[520] = 8'b10100110;
DRAM[521] = 8'b10100110;
DRAM[522] = 8'b10100110;
DRAM[523] = 8'b10100100;
DRAM[524] = 8'b10100011;
DRAM[525] = 8'b10011000;
DRAM[526] = 8'b10001010;
DRAM[527] = 8'b01110010;
DRAM[528] = 8'b01011010;
DRAM[529] = 8'b01011011;
DRAM[530] = 8'b01100010;
DRAM[531] = 8'b01100100;
DRAM[532] = 8'b01101010;
DRAM[533] = 8'b01101100;
DRAM[534] = 8'b01101001;
DRAM[535] = 8'b01101010;
DRAM[536] = 8'b01100110;
DRAM[537] = 8'b01100111;
DRAM[538] = 8'b01101111;
DRAM[539] = 8'b01110100;
DRAM[540] = 8'b01111001;
DRAM[541] = 8'b01111010;
DRAM[542] = 8'b01111010;
DRAM[543] = 8'b01111110;
DRAM[544] = 8'b10000001;
DRAM[545] = 8'b10000011;
DRAM[546] = 8'b10000010;
DRAM[547] = 8'b10000011;
DRAM[548] = 8'b10000100;
DRAM[549] = 8'b10000100;
DRAM[550] = 8'b10000011;
DRAM[551] = 8'b10000011;
DRAM[552] = 8'b10000100;
DRAM[553] = 8'b10000011;
DRAM[554] = 8'b10000101;
DRAM[555] = 8'b10000110;
DRAM[556] = 8'b10000101;
DRAM[557] = 8'b10000100;
DRAM[558] = 8'b10000011;
DRAM[559] = 8'b10000100;
DRAM[560] = 8'b10000011;
DRAM[561] = 8'b10001000;
DRAM[562] = 8'b10000100;
DRAM[563] = 8'b10000101;
DRAM[564] = 8'b10000101;
DRAM[565] = 8'b10000100;
DRAM[566] = 8'b10000100;
DRAM[567] = 8'b10000001;
DRAM[568] = 8'b10000001;
DRAM[569] = 8'b10000101;
DRAM[570] = 8'b10000001;
DRAM[571] = 8'b10000011;
DRAM[572] = 8'b10000110;
DRAM[573] = 8'b10001000;
DRAM[574] = 8'b10000100;
DRAM[575] = 8'b10000100;
DRAM[576] = 8'b10000110;
DRAM[577] = 8'b10000100;
DRAM[578] = 8'b10000001;
DRAM[579] = 8'b10000000;
DRAM[580] = 8'b10000011;
DRAM[581] = 8'b10000011;
DRAM[582] = 8'b01111101;
DRAM[583] = 8'b01111111;
DRAM[584] = 8'b10000000;
DRAM[585] = 8'b10000010;
DRAM[586] = 8'b01111110;
DRAM[587] = 8'b10000100;
DRAM[588] = 8'b01111011;
DRAM[589] = 8'b01111010;
DRAM[590] = 8'b01110011;
DRAM[591] = 8'b01110000;
DRAM[592] = 8'b01101011;
DRAM[593] = 8'b01100110;
DRAM[594] = 8'b01111000;
DRAM[595] = 8'b10001100;
DRAM[596] = 8'b10010110;
DRAM[597] = 8'b10011101;
DRAM[598] = 8'b10100010;
DRAM[599] = 8'b10100011;
DRAM[600] = 8'b10100001;
DRAM[601] = 8'b10100010;
DRAM[602] = 8'b10100011;
DRAM[603] = 8'b10100010;
DRAM[604] = 8'b10011110;
DRAM[605] = 8'b10011110;
DRAM[606] = 8'b10011101;
DRAM[607] = 8'b10011011;
DRAM[608] = 8'b10011010;
DRAM[609] = 8'b10011001;
DRAM[610] = 8'b10010111;
DRAM[611] = 8'b10010111;
DRAM[612] = 8'b10011000;
DRAM[613] = 8'b10010101;
DRAM[614] = 8'b10011111;
DRAM[615] = 8'b11001011;
DRAM[616] = 8'b11010111;
DRAM[617] = 8'b11011011;
DRAM[618] = 8'b11010100;
DRAM[619] = 8'b10011101;
DRAM[620] = 8'b01101000;
DRAM[621] = 8'b01101100;
DRAM[622] = 8'b01110100;
DRAM[623] = 8'b01110101;
DRAM[624] = 8'b01110111;
DRAM[625] = 8'b01111000;
DRAM[626] = 8'b01111100;
DRAM[627] = 8'b01111010;
DRAM[628] = 8'b01111100;
DRAM[629] = 8'b01111111;
DRAM[630] = 8'b01111101;
DRAM[631] = 8'b10000000;
DRAM[632] = 8'b10000010;
DRAM[633] = 8'b10000110;
DRAM[634] = 8'b01111110;
DRAM[635] = 8'b01001111;
DRAM[636] = 8'b00110000;
DRAM[637] = 8'b00101101;
DRAM[638] = 8'b00110000;
DRAM[639] = 8'b00101111;
DRAM[640] = 8'b10011010;
DRAM[641] = 8'b10011100;
DRAM[642] = 8'b10011110;
DRAM[643] = 8'b10011101;
DRAM[644] = 8'b10011100;
DRAM[645] = 8'b10011010;
DRAM[646] = 8'b10011100;
DRAM[647] = 8'b10100010;
DRAM[648] = 8'b10100110;
DRAM[649] = 8'b10100101;
DRAM[650] = 8'b10100100;
DRAM[651] = 8'b10100011;
DRAM[652] = 8'b10100010;
DRAM[653] = 8'b10011000;
DRAM[654] = 8'b10001001;
DRAM[655] = 8'b01110001;
DRAM[656] = 8'b01011010;
DRAM[657] = 8'b01011110;
DRAM[658] = 8'b01100001;
DRAM[659] = 8'b01101000;
DRAM[660] = 8'b01101000;
DRAM[661] = 8'b01101000;
DRAM[662] = 8'b01101000;
DRAM[663] = 8'b01100111;
DRAM[664] = 8'b01101000;
DRAM[665] = 8'b01101000;
DRAM[666] = 8'b01101101;
DRAM[667] = 8'b01110001;
DRAM[668] = 8'b01110110;
DRAM[669] = 8'b01111001;
DRAM[670] = 8'b01111110;
DRAM[671] = 8'b01111100;
DRAM[672] = 8'b10000001;
DRAM[673] = 8'b10000001;
DRAM[674] = 8'b10000001;
DRAM[675] = 8'b10000000;
DRAM[676] = 8'b10000101;
DRAM[677] = 8'b10000001;
DRAM[678] = 8'b10000001;
DRAM[679] = 8'b10000010;
DRAM[680] = 8'b10000011;
DRAM[681] = 8'b10000011;
DRAM[682] = 8'b10000011;
DRAM[683] = 8'b10000011;
DRAM[684] = 8'b10000010;
DRAM[685] = 8'b10000011;
DRAM[686] = 8'b10000010;
DRAM[687] = 8'b10000011;
DRAM[688] = 8'b10000011;
DRAM[689] = 8'b10000011;
DRAM[690] = 8'b10000000;
DRAM[691] = 8'b10000010;
DRAM[692] = 8'b01111111;
DRAM[693] = 8'b10000001;
DRAM[694] = 8'b10000010;
DRAM[695] = 8'b10000001;
DRAM[696] = 8'b10000001;
DRAM[697] = 8'b10000001;
DRAM[698] = 8'b10000000;
DRAM[699] = 8'b10000010;
DRAM[700] = 8'b10000100;
DRAM[701] = 8'b10000110;
DRAM[702] = 8'b10000111;
DRAM[703] = 8'b10000000;
DRAM[704] = 8'b10000011;
DRAM[705] = 8'b10000011;
DRAM[706] = 8'b10000011;
DRAM[707] = 8'b10000000;
DRAM[708] = 8'b10000000;
DRAM[709] = 8'b01111110;
DRAM[710] = 8'b01111110;
DRAM[711] = 8'b01111110;
DRAM[712] = 8'b10000000;
DRAM[713] = 8'b01111111;
DRAM[714] = 8'b01111111;
DRAM[715] = 8'b10000000;
DRAM[716] = 8'b01111101;
DRAM[717] = 8'b01111000;
DRAM[718] = 8'b01111000;
DRAM[719] = 8'b01110000;
DRAM[720] = 8'b01101100;
DRAM[721] = 8'b01101001;
DRAM[722] = 8'b01110001;
DRAM[723] = 8'b10000111;
DRAM[724] = 8'b10010110;
DRAM[725] = 8'b10011100;
DRAM[726] = 8'b10100011;
DRAM[727] = 8'b10100100;
DRAM[728] = 8'b10100001;
DRAM[729] = 8'b10100000;
DRAM[730] = 8'b10100001;
DRAM[731] = 8'b10100000;
DRAM[732] = 8'b10100000;
DRAM[733] = 8'b10011100;
DRAM[734] = 8'b10011100;
DRAM[735] = 8'b10011010;
DRAM[736] = 8'b10011000;
DRAM[737] = 8'b10010111;
DRAM[738] = 8'b10010111;
DRAM[739] = 8'b10010111;
DRAM[740] = 8'b10010110;
DRAM[741] = 8'b10010111;
DRAM[742] = 8'b10010010;
DRAM[743] = 8'b10110111;
DRAM[744] = 8'b11010001;
DRAM[745] = 8'b11011001;
DRAM[746] = 8'b11011011;
DRAM[747] = 8'b11000101;
DRAM[748] = 8'b01111001;
DRAM[749] = 8'b01101100;
DRAM[750] = 8'b01101110;
DRAM[751] = 8'b01110110;
DRAM[752] = 8'b01110100;
DRAM[753] = 8'b01111010;
DRAM[754] = 8'b01111010;
DRAM[755] = 8'b01111011;
DRAM[756] = 8'b01111011;
DRAM[757] = 8'b10000001;
DRAM[758] = 8'b01111111;
DRAM[759] = 8'b10000100;
DRAM[760] = 8'b10000111;
DRAM[761] = 8'b10000011;
DRAM[762] = 8'b01001001;
DRAM[763] = 8'b00110100;
DRAM[764] = 8'b00101111;
DRAM[765] = 8'b00110000;
DRAM[766] = 8'b00101110;
DRAM[767] = 8'b00110011;
DRAM[768] = 8'b10011011;
DRAM[769] = 8'b10011100;
DRAM[770] = 8'b10100000;
DRAM[771] = 8'b10011110;
DRAM[772] = 8'b10011110;
DRAM[773] = 8'b10011101;
DRAM[774] = 8'b10011110;
DRAM[775] = 8'b10100101;
DRAM[776] = 8'b10100110;
DRAM[777] = 8'b10100101;
DRAM[778] = 8'b10100011;
DRAM[779] = 8'b10011110;
DRAM[780] = 8'b10100000;
DRAM[781] = 8'b10011011;
DRAM[782] = 8'b10001001;
DRAM[783] = 8'b01101101;
DRAM[784] = 8'b01011001;
DRAM[785] = 8'b01011001;
DRAM[786] = 8'b01100000;
DRAM[787] = 8'b01100110;
DRAM[788] = 8'b01101010;
DRAM[789] = 8'b01101001;
DRAM[790] = 8'b01101010;
DRAM[791] = 8'b01100101;
DRAM[792] = 8'b01100100;
DRAM[793] = 8'b01101010;
DRAM[794] = 8'b01101100;
DRAM[795] = 8'b01110010;
DRAM[796] = 8'b01111000;
DRAM[797] = 8'b01111001;
DRAM[798] = 8'b01111101;
DRAM[799] = 8'b01111110;
DRAM[800] = 8'b01111111;
DRAM[801] = 8'b01111101;
DRAM[802] = 8'b01111111;
DRAM[803] = 8'b10000010;
DRAM[804] = 8'b10000000;
DRAM[805] = 8'b10000000;
DRAM[806] = 8'b10000010;
DRAM[807] = 8'b10000010;
DRAM[808] = 8'b10000010;
DRAM[809] = 8'b10000000;
DRAM[810] = 8'b10000010;
DRAM[811] = 8'b10000100;
DRAM[812] = 8'b10000001;
DRAM[813] = 8'b10000001;
DRAM[814] = 8'b10000001;
DRAM[815] = 8'b10000101;
DRAM[816] = 8'b10000110;
DRAM[817] = 8'b10000010;
DRAM[818] = 8'b01111110;
DRAM[819] = 8'b01111110;
DRAM[820] = 8'b01111011;
DRAM[821] = 8'b01111110;
DRAM[822] = 8'b01111111;
DRAM[823] = 8'b01111111;
DRAM[824] = 8'b01111111;
DRAM[825] = 8'b01111110;
DRAM[826] = 8'b01111110;
DRAM[827] = 8'b10000001;
DRAM[828] = 8'b10000000;
DRAM[829] = 8'b10000000;
DRAM[830] = 8'b10000100;
DRAM[831] = 8'b10000011;
DRAM[832] = 8'b10000011;
DRAM[833] = 8'b10000110;
DRAM[834] = 8'b10000001;
DRAM[835] = 8'b01111111;
DRAM[836] = 8'b10000000;
DRAM[837] = 8'b01111101;
DRAM[838] = 8'b01111101;
DRAM[839] = 8'b01111101;
DRAM[840] = 8'b10000000;
DRAM[841] = 8'b01111101;
DRAM[842] = 8'b01111111;
DRAM[843] = 8'b10000000;
DRAM[844] = 8'b01111100;
DRAM[845] = 8'b01111010;
DRAM[846] = 8'b01111011;
DRAM[847] = 8'b01110000;
DRAM[848] = 8'b01101100;
DRAM[849] = 8'b01101001;
DRAM[850] = 8'b01110101;
DRAM[851] = 8'b10000101;
DRAM[852] = 8'b10010101;
DRAM[853] = 8'b10011100;
DRAM[854] = 8'b10100010;
DRAM[855] = 8'b10100010;
DRAM[856] = 8'b10100100;
DRAM[857] = 8'b10100000;
DRAM[858] = 8'b10011111;
DRAM[859] = 8'b10011110;
DRAM[860] = 8'b10011111;
DRAM[861] = 8'b10011101;
DRAM[862] = 8'b10011011;
DRAM[863] = 8'b10011110;
DRAM[864] = 8'b10011011;
DRAM[865] = 8'b10011010;
DRAM[866] = 8'b10011000;
DRAM[867] = 8'b10010111;
DRAM[868] = 8'b10011000;
DRAM[869] = 8'b10010101;
DRAM[870] = 8'b10010100;
DRAM[871] = 8'b10011011;
DRAM[872] = 8'b11001001;
DRAM[873] = 8'b11010111;
DRAM[874] = 8'b11011011;
DRAM[875] = 8'b11011000;
DRAM[876] = 8'b10101100;
DRAM[877] = 8'b01101000;
DRAM[878] = 8'b01110000;
DRAM[879] = 8'b01110011;
DRAM[880] = 8'b01111010;
DRAM[881] = 8'b01111011;
DRAM[882] = 8'b01111100;
DRAM[883] = 8'b01111011;
DRAM[884] = 8'b01111001;
DRAM[885] = 8'b01111100;
DRAM[886] = 8'b10000000;
DRAM[887] = 8'b10000101;
DRAM[888] = 8'b10000010;
DRAM[889] = 8'b01001000;
DRAM[890] = 8'b00111010;
DRAM[891] = 8'b00101110;
DRAM[892] = 8'b00101100;
DRAM[893] = 8'b00101110;
DRAM[894] = 8'b00110010;
DRAM[895] = 8'b00110101;
DRAM[896] = 8'b10011110;
DRAM[897] = 8'b10011110;
DRAM[898] = 8'b10011110;
DRAM[899] = 8'b10011101;
DRAM[900] = 8'b10100001;
DRAM[901] = 8'b10100000;
DRAM[902] = 8'b10100110;
DRAM[903] = 8'b10101001;
DRAM[904] = 8'b10101001;
DRAM[905] = 8'b10100011;
DRAM[906] = 8'b10011110;
DRAM[907] = 8'b10011100;
DRAM[908] = 8'b10100100;
DRAM[909] = 8'b10011111;
DRAM[910] = 8'b10001001;
DRAM[911] = 8'b01101100;
DRAM[912] = 8'b01011010;
DRAM[913] = 8'b01011010;
DRAM[914] = 8'b01100101;
DRAM[915] = 8'b01101000;
DRAM[916] = 8'b01101010;
DRAM[917] = 8'b01101001;
DRAM[918] = 8'b01101010;
DRAM[919] = 8'b01101000;
DRAM[920] = 8'b01101000;
DRAM[921] = 8'b01101011;
DRAM[922] = 8'b01101110;
DRAM[923] = 8'b01110011;
DRAM[924] = 8'b01111000;
DRAM[925] = 8'b01111011;
DRAM[926] = 8'b01111010;
DRAM[927] = 8'b01111100;
DRAM[928] = 8'b10000001;
DRAM[929] = 8'b10000010;
DRAM[930] = 8'b01111101;
DRAM[931] = 8'b01111111;
DRAM[932] = 8'b01111110;
DRAM[933] = 8'b10000000;
DRAM[934] = 8'b10000001;
DRAM[935] = 8'b10000000;
DRAM[936] = 8'b10000011;
DRAM[937] = 8'b10000010;
DRAM[938] = 8'b10000001;
DRAM[939] = 8'b10000000;
DRAM[940] = 8'b10000000;
DRAM[941] = 8'b10000001;
DRAM[942] = 8'b10000000;
DRAM[943] = 8'b10000011;
DRAM[944] = 8'b10000101;
DRAM[945] = 8'b10000101;
DRAM[946] = 8'b01111111;
DRAM[947] = 8'b01111110;
DRAM[948] = 8'b01111001;
DRAM[949] = 8'b01111100;
DRAM[950] = 8'b01111100;
DRAM[951] = 8'b10000000;
DRAM[952] = 8'b01111100;
DRAM[953] = 8'b01111110;
DRAM[954] = 8'b01111011;
DRAM[955] = 8'b01111110;
DRAM[956] = 8'b10000001;
DRAM[957] = 8'b10000000;
DRAM[958] = 8'b01111111;
DRAM[959] = 8'b10000010;
DRAM[960] = 8'b10000011;
DRAM[961] = 8'b10000011;
DRAM[962] = 8'b01111101;
DRAM[963] = 8'b01111110;
DRAM[964] = 8'b10000000;
DRAM[965] = 8'b01111111;
DRAM[966] = 8'b01111110;
DRAM[967] = 8'b01111110;
DRAM[968] = 8'b01111110;
DRAM[969] = 8'b01111101;
DRAM[970] = 8'b01111101;
DRAM[971] = 8'b10000000;
DRAM[972] = 8'b01111101;
DRAM[973] = 8'b01110111;
DRAM[974] = 8'b01110110;
DRAM[975] = 8'b01110011;
DRAM[976] = 8'b01101110;
DRAM[977] = 8'b01101100;
DRAM[978] = 8'b01110100;
DRAM[979] = 8'b10000100;
DRAM[980] = 8'b10010000;
DRAM[981] = 8'b10011011;
DRAM[982] = 8'b10011100;
DRAM[983] = 8'b10100000;
DRAM[984] = 8'b10100001;
DRAM[985] = 8'b10011110;
DRAM[986] = 8'b10011110;
DRAM[987] = 8'b10011111;
DRAM[988] = 8'b10011101;
DRAM[989] = 8'b10011110;
DRAM[990] = 8'b10011100;
DRAM[991] = 8'b10011101;
DRAM[992] = 8'b10011010;
DRAM[993] = 8'b10011101;
DRAM[994] = 8'b10011100;
DRAM[995] = 8'b10011001;
DRAM[996] = 8'b10011010;
DRAM[997] = 8'b10010101;
DRAM[998] = 8'b10010010;
DRAM[999] = 8'b10001111;
DRAM[1000] = 8'b10101111;
DRAM[1001] = 8'b11010001;
DRAM[1002] = 8'b11011010;
DRAM[1003] = 8'b11011101;
DRAM[1004] = 8'b11010010;
DRAM[1005] = 8'b10000011;
DRAM[1006] = 8'b01101100;
DRAM[1007] = 8'b01110001;
DRAM[1008] = 8'b01110110;
DRAM[1009] = 8'b01111010;
DRAM[1010] = 8'b01111011;
DRAM[1011] = 8'b01111000;
DRAM[1012] = 8'b01111010;
DRAM[1013] = 8'b01111111;
DRAM[1014] = 8'b10000000;
DRAM[1015] = 8'b01111101;
DRAM[1016] = 8'b01001000;
DRAM[1017] = 8'b00101100;
DRAM[1018] = 8'b00101100;
DRAM[1019] = 8'b00110001;
DRAM[1020] = 8'b00110001;
DRAM[1021] = 8'b00110001;
DRAM[1022] = 8'b00101111;
DRAM[1023] = 8'b00110110;
DRAM[1024] = 8'b10011110;
DRAM[1025] = 8'b10011101;
DRAM[1026] = 8'b10100000;
DRAM[1027] = 8'b10100001;
DRAM[1028] = 8'b10100010;
DRAM[1029] = 8'b10100101;
DRAM[1030] = 8'b10100111;
DRAM[1031] = 8'b10101001;
DRAM[1032] = 8'b10101000;
DRAM[1033] = 8'b10100010;
DRAM[1034] = 8'b10011110;
DRAM[1035] = 8'b10011110;
DRAM[1036] = 8'b10100011;
DRAM[1037] = 8'b10011011;
DRAM[1038] = 8'b10001010;
DRAM[1039] = 8'b01101100;
DRAM[1040] = 8'b01011010;
DRAM[1041] = 8'b01011011;
DRAM[1042] = 8'b01100100;
DRAM[1043] = 8'b01101000;
DRAM[1044] = 8'b01101000;
DRAM[1045] = 8'b01101010;
DRAM[1046] = 8'b01101001;
DRAM[1047] = 8'b01100110;
DRAM[1048] = 8'b01100110;
DRAM[1049] = 8'b01101010;
DRAM[1050] = 8'b01101101;
DRAM[1051] = 8'b01110011;
DRAM[1052] = 8'b01110110;
DRAM[1053] = 8'b01111010;
DRAM[1054] = 8'b01111011;
DRAM[1055] = 8'b01111110;
DRAM[1056] = 8'b01111101;
DRAM[1057] = 8'b10000010;
DRAM[1058] = 8'b01111111;
DRAM[1059] = 8'b10000001;
DRAM[1060] = 8'b10000001;
DRAM[1061] = 8'b01111111;
DRAM[1062] = 8'b01111111;
DRAM[1063] = 8'b10000011;
DRAM[1064] = 8'b10000010;
DRAM[1065] = 8'b01111111;
DRAM[1066] = 8'b10000100;
DRAM[1067] = 8'b10000001;
DRAM[1068] = 8'b10000001;
DRAM[1069] = 8'b10000001;
DRAM[1070] = 8'b10000001;
DRAM[1071] = 8'b10000010;
DRAM[1072] = 8'b10000101;
DRAM[1073] = 8'b01111111;
DRAM[1074] = 8'b10000000;
DRAM[1075] = 8'b01111011;
DRAM[1076] = 8'b01111011;
DRAM[1077] = 8'b01111000;
DRAM[1078] = 8'b01111010;
DRAM[1079] = 8'b01111100;
DRAM[1080] = 8'b10000000;
DRAM[1081] = 8'b01111010;
DRAM[1082] = 8'b01111001;
DRAM[1083] = 8'b01111010;
DRAM[1084] = 8'b01111111;
DRAM[1085] = 8'b01111111;
DRAM[1086] = 8'b10000001;
DRAM[1087] = 8'b10000000;
DRAM[1088] = 8'b10000100;
DRAM[1089] = 8'b10000001;
DRAM[1090] = 8'b10000000;
DRAM[1091] = 8'b10000000;
DRAM[1092] = 8'b10000011;
DRAM[1093] = 8'b01111111;
DRAM[1094] = 8'b10000000;
DRAM[1095] = 8'b10000000;
DRAM[1096] = 8'b01111111;
DRAM[1097] = 8'b10000000;
DRAM[1098] = 8'b01111111;
DRAM[1099] = 8'b01111111;
DRAM[1100] = 8'b01111110;
DRAM[1101] = 8'b01111000;
DRAM[1102] = 8'b01110110;
DRAM[1103] = 8'b01101111;
DRAM[1104] = 8'b01110001;
DRAM[1105] = 8'b01101011;
DRAM[1106] = 8'b01110110;
DRAM[1107] = 8'b10000011;
DRAM[1108] = 8'b10001101;
DRAM[1109] = 8'b10010111;
DRAM[1110] = 8'b10011011;
DRAM[1111] = 8'b10100000;
DRAM[1112] = 8'b10011110;
DRAM[1113] = 8'b10011101;
DRAM[1114] = 8'b10011110;
DRAM[1115] = 8'b10011110;
DRAM[1116] = 8'b10011110;
DRAM[1117] = 8'b10011110;
DRAM[1118] = 8'b10011110;
DRAM[1119] = 8'b10011100;
DRAM[1120] = 8'b10011100;
DRAM[1121] = 8'b10011101;
DRAM[1122] = 8'b10011010;
DRAM[1123] = 8'b10011100;
DRAM[1124] = 8'b10011010;
DRAM[1125] = 8'b10010111;
DRAM[1126] = 8'b10010101;
DRAM[1127] = 8'b10010001;
DRAM[1128] = 8'b10010100;
DRAM[1129] = 8'b11000101;
DRAM[1130] = 8'b11011000;
DRAM[1131] = 8'b11011110;
DRAM[1132] = 8'b11011110;
DRAM[1133] = 8'b10111011;
DRAM[1134] = 8'b01110000;
DRAM[1135] = 8'b01101010;
DRAM[1136] = 8'b01110010;
DRAM[1137] = 8'b01110100;
DRAM[1138] = 8'b01111011;
DRAM[1139] = 8'b01111010;
DRAM[1140] = 8'b01111101;
DRAM[1141] = 8'b10000011;
DRAM[1142] = 8'b10000001;
DRAM[1143] = 8'b01000101;
DRAM[1144] = 8'b00101100;
DRAM[1145] = 8'b00101011;
DRAM[1146] = 8'b00110100;
DRAM[1147] = 8'b00110011;
DRAM[1148] = 8'b00110101;
DRAM[1149] = 8'b00110001;
DRAM[1150] = 8'b00110011;
DRAM[1151] = 8'b00110100;
DRAM[1152] = 8'b10100000;
DRAM[1153] = 8'b10011110;
DRAM[1154] = 8'b10100100;
DRAM[1155] = 8'b10100011;
DRAM[1156] = 8'b10100110;
DRAM[1157] = 8'b10101000;
DRAM[1158] = 8'b10100111;
DRAM[1159] = 8'b10100101;
DRAM[1160] = 8'b10100011;
DRAM[1161] = 8'b10100001;
DRAM[1162] = 8'b10011101;
DRAM[1163] = 8'b10100001;
DRAM[1164] = 8'b10100000;
DRAM[1165] = 8'b10011010;
DRAM[1166] = 8'b10001010;
DRAM[1167] = 8'b01101101;
DRAM[1168] = 8'b01010110;
DRAM[1169] = 8'b01010110;
DRAM[1170] = 8'b01100000;
DRAM[1171] = 8'b01100110;
DRAM[1172] = 8'b01101001;
DRAM[1173] = 8'b01100101;
DRAM[1174] = 8'b01101000;
DRAM[1175] = 8'b01101000;
DRAM[1176] = 8'b01101000;
DRAM[1177] = 8'b01101000;
DRAM[1178] = 8'b01101110;
DRAM[1179] = 8'b01110010;
DRAM[1180] = 8'b01110100;
DRAM[1181] = 8'b01111001;
DRAM[1182] = 8'b01110110;
DRAM[1183] = 8'b01111011;
DRAM[1184] = 8'b01111100;
DRAM[1185] = 8'b01111100;
DRAM[1186] = 8'b01111101;
DRAM[1187] = 8'b01111111;
DRAM[1188] = 8'b01111100;
DRAM[1189] = 8'b01111101;
DRAM[1190] = 8'b10000001;
DRAM[1191] = 8'b10000000;
DRAM[1192] = 8'b10000000;
DRAM[1193] = 8'b01111110;
DRAM[1194] = 8'b01111110;
DRAM[1195] = 8'b10000011;
DRAM[1196] = 8'b10000011;
DRAM[1197] = 8'b10000101;
DRAM[1198] = 8'b10000000;
DRAM[1199] = 8'b10000010;
DRAM[1200] = 8'b10000000;
DRAM[1201] = 8'b10000001;
DRAM[1202] = 8'b01111100;
DRAM[1203] = 8'b01111101;
DRAM[1204] = 8'b01111010;
DRAM[1205] = 8'b01111100;
DRAM[1206] = 8'b01111100;
DRAM[1207] = 8'b01111011;
DRAM[1208] = 8'b01111001;
DRAM[1209] = 8'b01110111;
DRAM[1210] = 8'b01111000;
DRAM[1211] = 8'b01111001;
DRAM[1212] = 8'b01111101;
DRAM[1213] = 8'b10000000;
DRAM[1214] = 8'b10000001;
DRAM[1215] = 8'b10000001;
DRAM[1216] = 8'b10000010;
DRAM[1217] = 8'b10000010;
DRAM[1218] = 8'b10000000;
DRAM[1219] = 8'b01111110;
DRAM[1220] = 8'b10000010;
DRAM[1221] = 8'b01111111;
DRAM[1222] = 8'b10000001;
DRAM[1223] = 8'b01111100;
DRAM[1224] = 8'b01111101;
DRAM[1225] = 8'b01111110;
DRAM[1226] = 8'b01111111;
DRAM[1227] = 8'b01111111;
DRAM[1228] = 8'b01111100;
DRAM[1229] = 8'b01111010;
DRAM[1230] = 8'b01110011;
DRAM[1231] = 8'b01110011;
DRAM[1232] = 8'b01110001;
DRAM[1233] = 8'b01101011;
DRAM[1234] = 8'b01110010;
DRAM[1235] = 8'b10000010;
DRAM[1236] = 8'b10001100;
DRAM[1237] = 8'b10010100;
DRAM[1238] = 8'b10011000;
DRAM[1239] = 8'b10011010;
DRAM[1240] = 8'b10011100;
DRAM[1241] = 8'b10011111;
DRAM[1242] = 8'b10011011;
DRAM[1243] = 8'b10011100;
DRAM[1244] = 8'b10011100;
DRAM[1245] = 8'b10011011;
DRAM[1246] = 8'b10011110;
DRAM[1247] = 8'b10011010;
DRAM[1248] = 8'b10011100;
DRAM[1249] = 8'b10011011;
DRAM[1250] = 8'b10011011;
DRAM[1251] = 8'b10011100;
DRAM[1252] = 8'b10011001;
DRAM[1253] = 8'b10010101;
DRAM[1254] = 8'b10010100;
DRAM[1255] = 8'b10010001;
DRAM[1256] = 8'b10001110;
DRAM[1257] = 8'b10100101;
DRAM[1258] = 8'b11010001;
DRAM[1259] = 8'b11011100;
DRAM[1260] = 8'b11011111;
DRAM[1261] = 8'b11011000;
DRAM[1262] = 8'b10011100;
DRAM[1263] = 8'b01100010;
DRAM[1264] = 8'b01101101;
DRAM[1265] = 8'b01110001;
DRAM[1266] = 8'b01111000;
DRAM[1267] = 8'b01111100;
DRAM[1268] = 8'b10000011;
DRAM[1269] = 8'b01111110;
DRAM[1270] = 8'b01000111;
DRAM[1271] = 8'b00101011;
DRAM[1272] = 8'b00101100;
DRAM[1273] = 8'b00101111;
DRAM[1274] = 8'b00111010;
DRAM[1275] = 8'b00111001;
DRAM[1276] = 8'b00111001;
DRAM[1277] = 8'b00110100;
DRAM[1278] = 8'b00101111;
DRAM[1279] = 8'b00110000;
DRAM[1280] = 8'b10100000;
DRAM[1281] = 8'b10100010;
DRAM[1282] = 8'b10100001;
DRAM[1283] = 8'b10100011;
DRAM[1284] = 8'b10101001;
DRAM[1285] = 8'b10100101;
DRAM[1286] = 8'b10100000;
DRAM[1287] = 8'b10100001;
DRAM[1288] = 8'b10011110;
DRAM[1289] = 8'b10100000;
DRAM[1290] = 8'b10011110;
DRAM[1291] = 8'b10011111;
DRAM[1292] = 8'b10100001;
DRAM[1293] = 8'b10011011;
DRAM[1294] = 8'b10000110;
DRAM[1295] = 8'b01101100;
DRAM[1296] = 8'b01010011;
DRAM[1297] = 8'b01011010;
DRAM[1298] = 8'b01100001;
DRAM[1299] = 8'b01100110;
DRAM[1300] = 8'b01100110;
DRAM[1301] = 8'b01101000;
DRAM[1302] = 8'b01100110;
DRAM[1303] = 8'b01101000;
DRAM[1304] = 8'b01100110;
DRAM[1305] = 8'b01101000;
DRAM[1306] = 8'b01101100;
DRAM[1307] = 8'b01110000;
DRAM[1308] = 8'b01111010;
DRAM[1309] = 8'b01111000;
DRAM[1310] = 8'b01111000;
DRAM[1311] = 8'b01111100;
DRAM[1312] = 8'b01111100;
DRAM[1313] = 8'b01111010;
DRAM[1314] = 8'b01111101;
DRAM[1315] = 8'b01111110;
DRAM[1316] = 8'b01111100;
DRAM[1317] = 8'b01111110;
DRAM[1318] = 8'b01111111;
DRAM[1319] = 8'b01111111;
DRAM[1320] = 8'b10000010;
DRAM[1321] = 8'b10000001;
DRAM[1322] = 8'b01111111;
DRAM[1323] = 8'b10000000;
DRAM[1324] = 8'b10000001;
DRAM[1325] = 8'b10000010;
DRAM[1326] = 8'b10000000;
DRAM[1327] = 8'b10000000;
DRAM[1328] = 8'b10000000;
DRAM[1329] = 8'b10000000;
DRAM[1330] = 8'b01111110;
DRAM[1331] = 8'b10000000;
DRAM[1332] = 8'b01111101;
DRAM[1333] = 8'b01111101;
DRAM[1334] = 8'b01111010;
DRAM[1335] = 8'b01111000;
DRAM[1336] = 8'b01110101;
DRAM[1337] = 8'b01110110;
DRAM[1338] = 8'b01110110;
DRAM[1339] = 8'b01110111;
DRAM[1340] = 8'b01110110;
DRAM[1341] = 8'b01111110;
DRAM[1342] = 8'b01111111;
DRAM[1343] = 8'b10000001;
DRAM[1344] = 8'b10000010;
DRAM[1345] = 8'b01111110;
DRAM[1346] = 8'b10000010;
DRAM[1347] = 8'b10000000;
DRAM[1348] = 8'b10000000;
DRAM[1349] = 8'b10000001;
DRAM[1350] = 8'b01111110;
DRAM[1351] = 8'b01111111;
DRAM[1352] = 8'b10000000;
DRAM[1353] = 8'b01111111;
DRAM[1354] = 8'b01111100;
DRAM[1355] = 8'b01111111;
DRAM[1356] = 8'b01111010;
DRAM[1357] = 8'b01111010;
DRAM[1358] = 8'b01110100;
DRAM[1359] = 8'b01110011;
DRAM[1360] = 8'b01110001;
DRAM[1361] = 8'b01101110;
DRAM[1362] = 8'b01110011;
DRAM[1363] = 8'b01111110;
DRAM[1364] = 8'b10001011;
DRAM[1365] = 8'b10010001;
DRAM[1366] = 8'b10010101;
DRAM[1367] = 8'b10011000;
DRAM[1368] = 8'b10011010;
DRAM[1369] = 8'b10011101;
DRAM[1370] = 8'b10011011;
DRAM[1371] = 8'b10011010;
DRAM[1372] = 8'b10011010;
DRAM[1373] = 8'b10011011;
DRAM[1374] = 8'b10011001;
DRAM[1375] = 8'b10011011;
DRAM[1376] = 8'b10011010;
DRAM[1377] = 8'b10011011;
DRAM[1378] = 8'b10011010;
DRAM[1379] = 8'b10011000;
DRAM[1380] = 8'b10010101;
DRAM[1381] = 8'b10010011;
DRAM[1382] = 8'b10010001;
DRAM[1383] = 8'b10001111;
DRAM[1384] = 8'b10001110;
DRAM[1385] = 8'b10001111;
DRAM[1386] = 8'b11000011;
DRAM[1387] = 8'b11011000;
DRAM[1388] = 8'b11011110;
DRAM[1389] = 8'b11011111;
DRAM[1390] = 8'b11000111;
DRAM[1391] = 8'b01110011;
DRAM[1392] = 8'b01101010;
DRAM[1393] = 8'b01110000;
DRAM[1394] = 8'b01110011;
DRAM[1395] = 8'b01111010;
DRAM[1396] = 8'b10000000;
DRAM[1397] = 8'b01001110;
DRAM[1398] = 8'b00101101;
DRAM[1399] = 8'b00101011;
DRAM[1400] = 8'b00101101;
DRAM[1401] = 8'b00110111;
DRAM[1402] = 8'b00111100;
DRAM[1403] = 8'b00110111;
DRAM[1404] = 8'b00110101;
DRAM[1405] = 8'b00110000;
DRAM[1406] = 8'b00101110;
DRAM[1407] = 8'b00101101;
DRAM[1408] = 8'b10100010;
DRAM[1409] = 8'b10100000;
DRAM[1410] = 8'b10100001;
DRAM[1411] = 8'b10100111;
DRAM[1412] = 8'b10100111;
DRAM[1413] = 8'b10011101;
DRAM[1414] = 8'b10011001;
DRAM[1415] = 8'b10011000;
DRAM[1416] = 8'b10011001;
DRAM[1417] = 8'b10100011;
DRAM[1418] = 8'b10100001;
DRAM[1419] = 8'b10100010;
DRAM[1420] = 8'b10100010;
DRAM[1421] = 8'b10011011;
DRAM[1422] = 8'b10001000;
DRAM[1423] = 8'b01101101;
DRAM[1424] = 8'b01010100;
DRAM[1425] = 8'b01011000;
DRAM[1426] = 8'b01100010;
DRAM[1427] = 8'b01100110;
DRAM[1428] = 8'b01100111;
DRAM[1429] = 8'b01101010;
DRAM[1430] = 8'b01100110;
DRAM[1431] = 8'b01100111;
DRAM[1432] = 8'b01100101;
DRAM[1433] = 8'b01101010;
DRAM[1434] = 8'b01101101;
DRAM[1435] = 8'b01110100;
DRAM[1436] = 8'b01110111;
DRAM[1437] = 8'b01111000;
DRAM[1438] = 8'b01111011;
DRAM[1439] = 8'b01111010;
DRAM[1440] = 8'b01111100;
DRAM[1441] = 8'b01111110;
DRAM[1442] = 8'b01111110;
DRAM[1443] = 8'b01111101;
DRAM[1444] = 8'b01111101;
DRAM[1445] = 8'b10000000;
DRAM[1446] = 8'b01111110;
DRAM[1447] = 8'b10000100;
DRAM[1448] = 8'b01111111;
DRAM[1449] = 8'b01111110;
DRAM[1450] = 8'b10000000;
DRAM[1451] = 8'b10000001;
DRAM[1452] = 8'b10000011;
DRAM[1453] = 8'b10000000;
DRAM[1454] = 8'b01111110;
DRAM[1455] = 8'b01111110;
DRAM[1456] = 8'b10000001;
DRAM[1457] = 8'b01111110;
DRAM[1458] = 8'b01111111;
DRAM[1459] = 8'b10000010;
DRAM[1460] = 8'b10001001;
DRAM[1461] = 8'b10000101;
DRAM[1462] = 8'b10010010;
DRAM[1463] = 8'b10100101;
DRAM[1464] = 8'b10100111;
DRAM[1465] = 8'b10100110;
DRAM[1466] = 8'b10100011;
DRAM[1467] = 8'b10010110;
DRAM[1468] = 8'b10001001;
DRAM[1469] = 8'b01110111;
DRAM[1470] = 8'b01110101;
DRAM[1471] = 8'b01110111;
DRAM[1472] = 8'b01111011;
DRAM[1473] = 8'b01111100;
DRAM[1474] = 8'b01111100;
DRAM[1475] = 8'b01111111;
DRAM[1476] = 8'b10000001;
DRAM[1477] = 8'b10000011;
DRAM[1478] = 8'b10000000;
DRAM[1479] = 8'b01111110;
DRAM[1480] = 8'b01111101;
DRAM[1481] = 8'b01111101;
DRAM[1482] = 8'b01111100;
DRAM[1483] = 8'b01111110;
DRAM[1484] = 8'b01111100;
DRAM[1485] = 8'b01111010;
DRAM[1486] = 8'b01110101;
DRAM[1487] = 8'b01110100;
DRAM[1488] = 8'b01101111;
DRAM[1489] = 8'b01101010;
DRAM[1490] = 8'b01110000;
DRAM[1491] = 8'b01111101;
DRAM[1492] = 8'b10001011;
DRAM[1493] = 8'b10010011;
DRAM[1494] = 8'b10010001;
DRAM[1495] = 8'b10010101;
DRAM[1496] = 8'b10010111;
DRAM[1497] = 8'b10011011;
DRAM[1498] = 8'b10011010;
DRAM[1499] = 8'b10011011;
DRAM[1500] = 8'b10011011;
DRAM[1501] = 8'b10011001;
DRAM[1502] = 8'b10011011;
DRAM[1503] = 8'b10011010;
DRAM[1504] = 8'b10011010;
DRAM[1505] = 8'b10011001;
DRAM[1506] = 8'b10011000;
DRAM[1507] = 8'b10010100;
DRAM[1508] = 8'b10010100;
DRAM[1509] = 8'b10010000;
DRAM[1510] = 8'b10010010;
DRAM[1511] = 8'b10001111;
DRAM[1512] = 8'b10001110;
DRAM[1513] = 8'b10001101;
DRAM[1514] = 8'b10100011;
DRAM[1515] = 8'b11010000;
DRAM[1516] = 8'b11011011;
DRAM[1517] = 8'b11011111;
DRAM[1518] = 8'b11011010;
DRAM[1519] = 8'b10100011;
DRAM[1520] = 8'b01101101;
DRAM[1521] = 8'b01101111;
DRAM[1522] = 8'b01110011;
DRAM[1523] = 8'b01111001;
DRAM[1524] = 8'b01001000;
DRAM[1525] = 8'b00101101;
DRAM[1526] = 8'b00101111;
DRAM[1527] = 8'b00101110;
DRAM[1528] = 8'b00110001;
DRAM[1529] = 8'b00111000;
DRAM[1530] = 8'b00111100;
DRAM[1531] = 8'b00110100;
DRAM[1532] = 8'b00110010;
DRAM[1533] = 8'b00101011;
DRAM[1534] = 8'b00101110;
DRAM[1535] = 8'b00101110;
DRAM[1536] = 8'b10100001;
DRAM[1537] = 8'b10011111;
DRAM[1538] = 8'b10100010;
DRAM[1539] = 8'b10101010;
DRAM[1540] = 8'b10100100;
DRAM[1541] = 8'b10010110;
DRAM[1542] = 8'b10010001;
DRAM[1543] = 8'b10010000;
DRAM[1544] = 8'b10011001;
DRAM[1545] = 8'b10100011;
DRAM[1546] = 8'b10100000;
DRAM[1547] = 8'b10100000;
DRAM[1548] = 8'b10100011;
DRAM[1549] = 8'b10011011;
DRAM[1550] = 8'b10001010;
DRAM[1551] = 8'b01101110;
DRAM[1552] = 8'b01010110;
DRAM[1553] = 8'b01011000;
DRAM[1554] = 8'b01100000;
DRAM[1555] = 8'b01100011;
DRAM[1556] = 8'b01101000;
DRAM[1557] = 8'b01101000;
DRAM[1558] = 8'b01100110;
DRAM[1559] = 8'b01101000;
DRAM[1560] = 8'b01100111;
DRAM[1561] = 8'b01101100;
DRAM[1562] = 8'b01110000;
DRAM[1563] = 8'b01110010;
DRAM[1564] = 8'b01111000;
DRAM[1565] = 8'b01111000;
DRAM[1566] = 8'b01111000;
DRAM[1567] = 8'b01111101;
DRAM[1568] = 8'b01111101;
DRAM[1569] = 8'b01111111;
DRAM[1570] = 8'b01111101;
DRAM[1571] = 8'b01111110;
DRAM[1572] = 8'b10000001;
DRAM[1573] = 8'b10000000;
DRAM[1574] = 8'b10000010;
DRAM[1575] = 8'b10000000;
DRAM[1576] = 8'b10000001;
DRAM[1577] = 8'b10000000;
DRAM[1578] = 8'b10000000;
DRAM[1579] = 8'b10000010;
DRAM[1580] = 8'b10000010;
DRAM[1581] = 8'b01111111;
DRAM[1582] = 8'b10000000;
DRAM[1583] = 8'b01111101;
DRAM[1584] = 8'b10001010;
DRAM[1585] = 8'b10010011;
DRAM[1586] = 8'b10010100;
DRAM[1587] = 8'b10010011;
DRAM[1588] = 8'b10010100;
DRAM[1589] = 8'b10100011;
DRAM[1590] = 8'b10100011;
DRAM[1591] = 8'b10101010;
DRAM[1592] = 8'b10110100;
DRAM[1593] = 8'b10110011;
DRAM[1594] = 8'b10110101;
DRAM[1595] = 8'b10110011;
DRAM[1596] = 8'b10110110;
DRAM[1597] = 8'b10111100;
DRAM[1598] = 8'b10100100;
DRAM[1599] = 8'b10001100;
DRAM[1600] = 8'b01110111;
DRAM[1601] = 8'b01110110;
DRAM[1602] = 8'b01111010;
DRAM[1603] = 8'b01111011;
DRAM[1604] = 8'b10000000;
DRAM[1605] = 8'b10000011;
DRAM[1606] = 8'b10000000;
DRAM[1607] = 8'b01111100;
DRAM[1608] = 8'b01111111;
DRAM[1609] = 8'b01111111;
DRAM[1610] = 8'b01111111;
DRAM[1611] = 8'b01111110;
DRAM[1612] = 8'b01111001;
DRAM[1613] = 8'b01110110;
DRAM[1614] = 8'b01110110;
DRAM[1615] = 8'b01110000;
DRAM[1616] = 8'b01101111;
DRAM[1617] = 8'b01101010;
DRAM[1618] = 8'b01101101;
DRAM[1619] = 8'b01111101;
DRAM[1620] = 8'b10001001;
DRAM[1621] = 8'b10010000;
DRAM[1622] = 8'b10001111;
DRAM[1623] = 8'b10010011;
DRAM[1624] = 8'b10010100;
DRAM[1625] = 8'b10011000;
DRAM[1626] = 8'b10011010;
DRAM[1627] = 8'b10011011;
DRAM[1628] = 8'b10011000;
DRAM[1629] = 8'b10011001;
DRAM[1630] = 8'b10011000;
DRAM[1631] = 8'b10011010;
DRAM[1632] = 8'b10011000;
DRAM[1633] = 8'b10011000;
DRAM[1634] = 8'b10010101;
DRAM[1635] = 8'b10010010;
DRAM[1636] = 8'b10010000;
DRAM[1637] = 8'b10001111;
DRAM[1638] = 8'b10001110;
DRAM[1639] = 8'b10001110;
DRAM[1640] = 8'b10001101;
DRAM[1641] = 8'b10001101;
DRAM[1642] = 8'b10010001;
DRAM[1643] = 8'b10111000;
DRAM[1644] = 8'b11010110;
DRAM[1645] = 8'b11011101;
DRAM[1646] = 8'b11100000;
DRAM[1647] = 8'b11010000;
DRAM[1648] = 8'b10000100;
DRAM[1649] = 8'b01110010;
DRAM[1650] = 8'b01110100;
DRAM[1651] = 8'b01001100;
DRAM[1652] = 8'b00101010;
DRAM[1653] = 8'b00101011;
DRAM[1654] = 8'b00101011;
DRAM[1655] = 8'b00101111;
DRAM[1656] = 8'b00110101;
DRAM[1657] = 8'b00111001;
DRAM[1658] = 8'b00111000;
DRAM[1659] = 8'b00111000;
DRAM[1660] = 8'b00101011;
DRAM[1661] = 8'b00101100;
DRAM[1662] = 8'b00110000;
DRAM[1663] = 8'b00101100;
DRAM[1664] = 8'b10100000;
DRAM[1665] = 8'b10100011;
DRAM[1666] = 8'b10100111;
DRAM[1667] = 8'b10100101;
DRAM[1668] = 8'b10011100;
DRAM[1669] = 8'b10001110;
DRAM[1670] = 8'b10000101;
DRAM[1671] = 8'b10001100;
DRAM[1672] = 8'b10011100;
DRAM[1673] = 8'b10100100;
DRAM[1674] = 8'b10100010;
DRAM[1675] = 8'b10100011;
DRAM[1676] = 8'b10100101;
DRAM[1677] = 8'b10011100;
DRAM[1678] = 8'b10001001;
DRAM[1679] = 8'b01101101;
DRAM[1680] = 8'b01010001;
DRAM[1681] = 8'b01011000;
DRAM[1682] = 8'b01011100;
DRAM[1683] = 8'b01100001;
DRAM[1684] = 8'b01101010;
DRAM[1685] = 8'b01100110;
DRAM[1686] = 8'b01100111;
DRAM[1687] = 8'b01100111;
DRAM[1688] = 8'b01101001;
DRAM[1689] = 8'b01101100;
DRAM[1690] = 8'b01110001;
DRAM[1691] = 8'b01110100;
DRAM[1692] = 8'b01110111;
DRAM[1693] = 8'b01111000;
DRAM[1694] = 8'b01111001;
DRAM[1695] = 8'b01111101;
DRAM[1696] = 8'b01111101;
DRAM[1697] = 8'b01111101;
DRAM[1698] = 8'b01111100;
DRAM[1699] = 8'b10000001;
DRAM[1700] = 8'b10000011;
DRAM[1701] = 8'b01111110;
DRAM[1702] = 8'b01111111;
DRAM[1703] = 8'b10000000;
DRAM[1704] = 8'b01111111;
DRAM[1705] = 8'b01111111;
DRAM[1706] = 8'b10000001;
DRAM[1707] = 8'b10000000;
DRAM[1708] = 8'b10000000;
DRAM[1709] = 8'b10000000;
DRAM[1710] = 8'b10000000;
DRAM[1711] = 8'b10010010;
DRAM[1712] = 8'b10010001;
DRAM[1713] = 8'b10010110;
DRAM[1714] = 8'b10010000;
DRAM[1715] = 8'b10010100;
DRAM[1716] = 8'b10011001;
DRAM[1717] = 8'b10100101;
DRAM[1718] = 8'b10100011;
DRAM[1719] = 8'b10101011;
DRAM[1720] = 8'b10110011;
DRAM[1721] = 8'b10110001;
DRAM[1722] = 8'b10101110;
DRAM[1723] = 8'b10101100;
DRAM[1724] = 8'b10110010;
DRAM[1725] = 8'b10111001;
DRAM[1726] = 8'b10111010;
DRAM[1727] = 8'b11000010;
DRAM[1728] = 8'b10111001;
DRAM[1729] = 8'b10010100;
DRAM[1730] = 8'b01110001;
DRAM[1731] = 8'b01111100;
DRAM[1732] = 8'b01111010;
DRAM[1733] = 8'b01111110;
DRAM[1734] = 8'b01111110;
DRAM[1735] = 8'b10000000;
DRAM[1736] = 8'b01111100;
DRAM[1737] = 8'b01111110;
DRAM[1738] = 8'b01111010;
DRAM[1739] = 8'b01111100;
DRAM[1740] = 8'b01111001;
DRAM[1741] = 8'b01111000;
DRAM[1742] = 8'b01110000;
DRAM[1743] = 8'b01110010;
DRAM[1744] = 8'b01110001;
DRAM[1745] = 8'b01101001;
DRAM[1746] = 8'b01110011;
DRAM[1747] = 8'b10000000;
DRAM[1748] = 8'b10001011;
DRAM[1749] = 8'b10010010;
DRAM[1750] = 8'b10010000;
DRAM[1751] = 8'b10010000;
DRAM[1752] = 8'b10010011;
DRAM[1753] = 8'b10010110;
DRAM[1754] = 8'b10011001;
DRAM[1755] = 8'b10011001;
DRAM[1756] = 8'b10011011;
DRAM[1757] = 8'b10010111;
DRAM[1758] = 8'b10010110;
DRAM[1759] = 8'b10010101;
DRAM[1760] = 8'b10010100;
DRAM[1761] = 8'b10010011;
DRAM[1762] = 8'b10010001;
DRAM[1763] = 8'b10010000;
DRAM[1764] = 8'b10010000;
DRAM[1765] = 8'b10001100;
DRAM[1766] = 8'b10001101;
DRAM[1767] = 8'b10001011;
DRAM[1768] = 8'b10001110;
DRAM[1769] = 8'b10001101;
DRAM[1770] = 8'b10001101;
DRAM[1771] = 8'b10010101;
DRAM[1772] = 8'b11001011;
DRAM[1773] = 8'b11011011;
DRAM[1774] = 8'b11100000;
DRAM[1775] = 8'b11100000;
DRAM[1776] = 8'b10111110;
DRAM[1777] = 8'b01111000;
DRAM[1778] = 8'b01010101;
DRAM[1779] = 8'b00101110;
DRAM[1780] = 8'b00101010;
DRAM[1781] = 8'b00101110;
DRAM[1782] = 8'b00110001;
DRAM[1783] = 8'b00110100;
DRAM[1784] = 8'b00110110;
DRAM[1785] = 8'b00110100;
DRAM[1786] = 8'b00110011;
DRAM[1787] = 8'b00110000;
DRAM[1788] = 8'b00110100;
DRAM[1789] = 8'b00110000;
DRAM[1790] = 8'b00101111;
DRAM[1791] = 8'b00101101;
DRAM[1792] = 8'b10100000;
DRAM[1793] = 8'b10100111;
DRAM[1794] = 8'b10101100;
DRAM[1795] = 8'b10011110;
DRAM[1796] = 8'b10010011;
DRAM[1797] = 8'b01111110;
DRAM[1798] = 8'b01111010;
DRAM[1799] = 8'b10001110;
DRAM[1800] = 8'b10011110;
DRAM[1801] = 8'b10100101;
DRAM[1802] = 8'b10100101;
DRAM[1803] = 8'b10100100;
DRAM[1804] = 8'b10100011;
DRAM[1805] = 8'b10011011;
DRAM[1806] = 8'b10001101;
DRAM[1807] = 8'b01101011;
DRAM[1808] = 8'b01010010;
DRAM[1809] = 8'b01010011;
DRAM[1810] = 8'b01100001;
DRAM[1811] = 8'b01100001;
DRAM[1812] = 8'b01100000;
DRAM[1813] = 8'b01100101;
DRAM[1814] = 8'b01100011;
DRAM[1815] = 8'b01100100;
DRAM[1816] = 8'b01101010;
DRAM[1817] = 8'b01101001;
DRAM[1818] = 8'b01110000;
DRAM[1819] = 8'b01110001;
DRAM[1820] = 8'b01110101;
DRAM[1821] = 8'b01110111;
DRAM[1822] = 8'b01111010;
DRAM[1823] = 8'b01111001;
DRAM[1824] = 8'b01111100;
DRAM[1825] = 8'b01111001;
DRAM[1826] = 8'b01111010;
DRAM[1827] = 8'b01111110;
DRAM[1828] = 8'b01111111;
DRAM[1829] = 8'b01111111;
DRAM[1830] = 8'b01111111;
DRAM[1831] = 8'b01111110;
DRAM[1832] = 8'b01111110;
DRAM[1833] = 8'b10000000;
DRAM[1834] = 8'b10001111;
DRAM[1835] = 8'b10010000;
DRAM[1836] = 8'b10000111;
DRAM[1837] = 8'b01111010;
DRAM[1838] = 8'b10001000;
DRAM[1839] = 8'b10001011;
DRAM[1840] = 8'b10001111;
DRAM[1841] = 8'b10001010;
DRAM[1842] = 8'b10010001;
DRAM[1843] = 8'b10010111;
DRAM[1844] = 8'b10010010;
DRAM[1845] = 8'b10011101;
DRAM[1846] = 8'b10011111;
DRAM[1847] = 8'b10100101;
DRAM[1848] = 8'b10101010;
DRAM[1849] = 8'b10101100;
DRAM[1850] = 8'b10101111;
DRAM[1851] = 8'b10110010;
DRAM[1852] = 8'b10110001;
DRAM[1853] = 8'b10111001;
DRAM[1854] = 8'b10111010;
DRAM[1855] = 8'b10111110;
DRAM[1856] = 8'b11000100;
DRAM[1857] = 8'b11000011;
DRAM[1858] = 8'b10110000;
DRAM[1859] = 8'b01111000;
DRAM[1860] = 8'b01110100;
DRAM[1861] = 8'b01111001;
DRAM[1862] = 8'b01111100;
DRAM[1863] = 8'b01111100;
DRAM[1864] = 8'b01111010;
DRAM[1865] = 8'b01111101;
DRAM[1866] = 8'b01111101;
DRAM[1867] = 8'b01111010;
DRAM[1868] = 8'b01110011;
DRAM[1869] = 8'b01110101;
DRAM[1870] = 8'b01110001;
DRAM[1871] = 8'b01101111;
DRAM[1872] = 8'b01101110;
DRAM[1873] = 8'b01101010;
DRAM[1874] = 8'b01110000;
DRAM[1875] = 8'b01111100;
DRAM[1876] = 8'b10001011;
DRAM[1877] = 8'b10010000;
DRAM[1878] = 8'b10010011;
DRAM[1879] = 8'b10010001;
DRAM[1880] = 8'b10010010;
DRAM[1881] = 8'b10010100;
DRAM[1882] = 8'b10010110;
DRAM[1883] = 8'b10011000;
DRAM[1884] = 8'b10010110;
DRAM[1885] = 8'b10010100;
DRAM[1886] = 8'b10010001;
DRAM[1887] = 8'b10010010;
DRAM[1888] = 8'b10010001;
DRAM[1889] = 8'b10010000;
DRAM[1890] = 8'b10010010;
DRAM[1891] = 8'b10001110;
DRAM[1892] = 8'b10001101;
DRAM[1893] = 8'b10001100;
DRAM[1894] = 8'b10001011;
DRAM[1895] = 8'b10001011;
DRAM[1896] = 8'b10001011;
DRAM[1897] = 8'b10001101;
DRAM[1898] = 8'b10010000;
DRAM[1899] = 8'b10001010;
DRAM[1900] = 8'b10101100;
DRAM[1901] = 8'b11010101;
DRAM[1902] = 8'b11011111;
DRAM[1903] = 8'b11100011;
DRAM[1904] = 8'b11011101;
DRAM[1905] = 8'b10000000;
DRAM[1906] = 8'b00101100;
DRAM[1907] = 8'b00101001;
DRAM[1908] = 8'b00101110;
DRAM[1909] = 8'b00110000;
DRAM[1910] = 8'b00110111;
DRAM[1911] = 8'b00110110;
DRAM[1912] = 8'b00110100;
DRAM[1913] = 8'b00110001;
DRAM[1914] = 8'b00101111;
DRAM[1915] = 8'b00110010;
DRAM[1916] = 8'b00110011;
DRAM[1917] = 8'b00101110;
DRAM[1918] = 8'b00101100;
DRAM[1919] = 8'b00110001;
DRAM[1920] = 8'b10100011;
DRAM[1921] = 8'b10101011;
DRAM[1922] = 8'b10101000;
DRAM[1923] = 8'b10011011;
DRAM[1924] = 8'b10001001;
DRAM[1925] = 8'b01101001;
DRAM[1926] = 8'b01101111;
DRAM[1927] = 8'b10001101;
DRAM[1928] = 8'b10011100;
DRAM[1929] = 8'b10100111;
DRAM[1930] = 8'b10100101;
DRAM[1931] = 8'b10100110;
DRAM[1932] = 8'b10100101;
DRAM[1933] = 8'b10011101;
DRAM[1934] = 8'b10001111;
DRAM[1935] = 8'b01101100;
DRAM[1936] = 8'b01010010;
DRAM[1937] = 8'b01010000;
DRAM[1938] = 8'b01010100;
DRAM[1939] = 8'b01011110;
DRAM[1940] = 8'b01100011;
DRAM[1941] = 8'b01100001;
DRAM[1942] = 8'b01100010;
DRAM[1943] = 8'b01100110;
DRAM[1944] = 8'b01101000;
DRAM[1945] = 8'b01100111;
DRAM[1946] = 8'b01101100;
DRAM[1947] = 8'b01110000;
DRAM[1948] = 8'b01110100;
DRAM[1949] = 8'b01110110;
DRAM[1950] = 8'b01111011;
DRAM[1951] = 8'b01111001;
DRAM[1952] = 8'b01111100;
DRAM[1953] = 8'b01111010;
DRAM[1954] = 8'b01111010;
DRAM[1955] = 8'b01111111;
DRAM[1956] = 8'b01111110;
DRAM[1957] = 8'b01111101;
DRAM[1958] = 8'b01111110;
DRAM[1959] = 8'b10001110;
DRAM[1960] = 8'b10000000;
DRAM[1961] = 8'b10010010;
DRAM[1962] = 8'b10001000;
DRAM[1963] = 8'b10000010;
DRAM[1964] = 8'b01111100;
DRAM[1965] = 8'b01111011;
DRAM[1966] = 8'b10000001;
DRAM[1967] = 8'b10000111;
DRAM[1968] = 8'b10000011;
DRAM[1969] = 8'b10000101;
DRAM[1970] = 8'b10001001;
DRAM[1971] = 8'b10001101;
DRAM[1972] = 8'b10010100;
DRAM[1973] = 8'b10011001;
DRAM[1974] = 8'b10100010;
DRAM[1975] = 8'b10011100;
DRAM[1976] = 8'b10101101;
DRAM[1977] = 8'b10101010;
DRAM[1978] = 8'b10110011;
DRAM[1979] = 8'b10110100;
DRAM[1980] = 8'b10111001;
DRAM[1981] = 8'b10110110;
DRAM[1982] = 8'b10111100;
DRAM[1983] = 8'b10111101;
DRAM[1984] = 8'b11000000;
DRAM[1985] = 8'b11000001;
DRAM[1986] = 8'b11000111;
DRAM[1987] = 8'b11000101;
DRAM[1988] = 8'b10010001;
DRAM[1989] = 8'b01110000;
DRAM[1990] = 8'b01110001;
DRAM[1991] = 8'b01110110;
DRAM[1992] = 8'b01110110;
DRAM[1993] = 8'b01111010;
DRAM[1994] = 8'b01111000;
DRAM[1995] = 8'b01111011;
DRAM[1996] = 8'b01110110;
DRAM[1997] = 8'b01110011;
DRAM[1998] = 8'b01110000;
DRAM[1999] = 8'b01101110;
DRAM[2000] = 8'b01101010;
DRAM[2001] = 8'b01100110;
DRAM[2002] = 8'b01101101;
DRAM[2003] = 8'b01111101;
DRAM[2004] = 8'b10001100;
DRAM[2005] = 8'b10010011;
DRAM[2006] = 8'b10010010;
DRAM[2007] = 8'b10010001;
DRAM[2008] = 8'b10010001;
DRAM[2009] = 8'b10010100;
DRAM[2010] = 8'b10010001;
DRAM[2011] = 8'b10010110;
DRAM[2012] = 8'b10010110;
DRAM[2013] = 8'b10010111;
DRAM[2014] = 8'b10010001;
DRAM[2015] = 8'b10001111;
DRAM[2016] = 8'b10001101;
DRAM[2017] = 8'b10010000;
DRAM[2018] = 8'b10010000;
DRAM[2019] = 8'b10010001;
DRAM[2020] = 8'b10001111;
DRAM[2021] = 8'b10001110;
DRAM[2022] = 8'b10001101;
DRAM[2023] = 8'b10001110;
DRAM[2024] = 8'b10001100;
DRAM[2025] = 8'b10001111;
DRAM[2026] = 8'b10001110;
DRAM[2027] = 8'b10001011;
DRAM[2028] = 8'b10001101;
DRAM[2029] = 8'b11000100;
DRAM[2030] = 8'b11011011;
DRAM[2031] = 8'b11100100;
DRAM[2032] = 8'b11011111;
DRAM[2033] = 8'b01011001;
DRAM[2034] = 8'b00100111;
DRAM[2035] = 8'b00101100;
DRAM[2036] = 8'b00101101;
DRAM[2037] = 8'b00110001;
DRAM[2038] = 8'b00111000;
DRAM[2039] = 8'b00110111;
DRAM[2040] = 8'b00110110;
DRAM[2041] = 8'b00101101;
DRAM[2042] = 8'b00101110;
DRAM[2043] = 8'b00110011;
DRAM[2044] = 8'b00101101;
DRAM[2045] = 8'b00101111;
DRAM[2046] = 8'b00101111;
DRAM[2047] = 8'b00110110;
DRAM[2048] = 8'b10101010;
DRAM[2049] = 8'b10101101;
DRAM[2050] = 8'b10100000;
DRAM[2051] = 8'b10010001;
DRAM[2052] = 8'b01110101;
DRAM[2053] = 8'b01010101;
DRAM[2054] = 8'b01101111;
DRAM[2055] = 8'b10001111;
DRAM[2056] = 8'b10100000;
DRAM[2057] = 8'b10100100;
DRAM[2058] = 8'b10100110;
DRAM[2059] = 8'b10100101;
DRAM[2060] = 8'b10100011;
DRAM[2061] = 8'b10011011;
DRAM[2062] = 8'b10001010;
DRAM[2063] = 8'b01101011;
DRAM[2064] = 8'b01001101;
DRAM[2065] = 8'b01010000;
DRAM[2066] = 8'b01010110;
DRAM[2067] = 8'b01011110;
DRAM[2068] = 8'b01011110;
DRAM[2069] = 8'b01100010;
DRAM[2070] = 8'b01100010;
DRAM[2071] = 8'b01100010;
DRAM[2072] = 8'b01100101;
DRAM[2073] = 8'b01101000;
DRAM[2074] = 8'b01101001;
DRAM[2075] = 8'b01101110;
DRAM[2076] = 8'b01110100;
DRAM[2077] = 8'b01110011;
DRAM[2078] = 8'b01110100;
DRAM[2079] = 8'b01110110;
DRAM[2080] = 8'b01111101;
DRAM[2081] = 8'b01111011;
DRAM[2082] = 8'b01111010;
DRAM[2083] = 8'b01111101;
DRAM[2084] = 8'b01111011;
DRAM[2085] = 8'b01111011;
DRAM[2086] = 8'b01111001;
DRAM[2087] = 8'b10010011;
DRAM[2088] = 8'b01101100;
DRAM[2089] = 8'b01111000;
DRAM[2090] = 8'b01111001;
DRAM[2091] = 8'b01110111;
DRAM[2092] = 8'b01111001;
DRAM[2093] = 8'b01111000;
DRAM[2094] = 8'b10000000;
DRAM[2095] = 8'b10000100;
DRAM[2096] = 8'b01111100;
DRAM[2097] = 8'b10000011;
DRAM[2098] = 8'b10001001;
DRAM[2099] = 8'b10001101;
DRAM[2100] = 8'b10001110;
DRAM[2101] = 8'b10010100;
DRAM[2102] = 8'b10011000;
DRAM[2103] = 8'b10011110;
DRAM[2104] = 8'b10101000;
DRAM[2105] = 8'b10101111;
DRAM[2106] = 8'b10110010;
DRAM[2107] = 8'b10110111;
DRAM[2108] = 8'b10111001;
DRAM[2109] = 8'b10111001;
DRAM[2110] = 8'b10111100;
DRAM[2111] = 8'b10111101;
DRAM[2112] = 8'b10111100;
DRAM[2113] = 8'b11000010;
DRAM[2114] = 8'b11000010;
DRAM[2115] = 8'b11000101;
DRAM[2116] = 8'b11000001;
DRAM[2117] = 8'b10101111;
DRAM[2118] = 8'b01110001;
DRAM[2119] = 8'b01101010;
DRAM[2120] = 8'b01110101;
DRAM[2121] = 8'b01110010;
DRAM[2122] = 8'b01110100;
DRAM[2123] = 8'b01110101;
DRAM[2124] = 8'b01110110;
DRAM[2125] = 8'b01110010;
DRAM[2126] = 8'b01110001;
DRAM[2127] = 8'b01101111;
DRAM[2128] = 8'b01101011;
DRAM[2129] = 8'b01101000;
DRAM[2130] = 8'b01101100;
DRAM[2131] = 8'b01111111;
DRAM[2132] = 8'b10001101;
DRAM[2133] = 8'b10010100;
DRAM[2134] = 8'b10010101;
DRAM[2135] = 8'b10010001;
DRAM[2136] = 8'b10010001;
DRAM[2137] = 8'b10001111;
DRAM[2138] = 8'b10001111;
DRAM[2139] = 8'b10001101;
DRAM[2140] = 8'b10010011;
DRAM[2141] = 8'b10010101;
DRAM[2142] = 8'b10010000;
DRAM[2143] = 8'b10001101;
DRAM[2144] = 8'b10001101;
DRAM[2145] = 8'b10001110;
DRAM[2146] = 8'b10010001;
DRAM[2147] = 8'b10001110;
DRAM[2148] = 8'b10001110;
DRAM[2149] = 8'b10001110;
DRAM[2150] = 8'b10001100;
DRAM[2151] = 8'b10001110;
DRAM[2152] = 8'b10001110;
DRAM[2153] = 8'b10010000;
DRAM[2154] = 8'b10001101;
DRAM[2155] = 8'b10001110;
DRAM[2156] = 8'b10001101;
DRAM[2157] = 8'b10011110;
DRAM[2158] = 8'b11011000;
DRAM[2159] = 8'b11011110;
DRAM[2160] = 8'b10001010;
DRAM[2161] = 8'b00100100;
DRAM[2162] = 8'b00101010;
DRAM[2163] = 8'b00101100;
DRAM[2164] = 8'b00110010;
DRAM[2165] = 8'b00111001;
DRAM[2166] = 8'b00110111;
DRAM[2167] = 8'b00111000;
DRAM[2168] = 8'b00101011;
DRAM[2169] = 8'b00101101;
DRAM[2170] = 8'b00110110;
DRAM[2171] = 8'b00110000;
DRAM[2172] = 8'b00101111;
DRAM[2173] = 8'b00110010;
DRAM[2174] = 8'b00110001;
DRAM[2175] = 8'b00100100;
DRAM[2176] = 8'b10101101;
DRAM[2177] = 8'b10100110;
DRAM[2178] = 8'b10011001;
DRAM[2179] = 8'b10000010;
DRAM[2180] = 8'b01011001;
DRAM[2181] = 8'b01001111;
DRAM[2182] = 8'b01101110;
DRAM[2183] = 8'b10001001;
DRAM[2184] = 8'b10011111;
DRAM[2185] = 8'b10101001;
DRAM[2186] = 8'b10100101;
DRAM[2187] = 8'b10100100;
DRAM[2188] = 8'b10100011;
DRAM[2189] = 8'b10011010;
DRAM[2190] = 8'b10000111;
DRAM[2191] = 8'b01101001;
DRAM[2192] = 8'b01001110;
DRAM[2193] = 8'b01010010;
DRAM[2194] = 8'b01010110;
DRAM[2195] = 8'b01011110;
DRAM[2196] = 8'b01100011;
DRAM[2197] = 8'b01100110;
DRAM[2198] = 8'b01100100;
DRAM[2199] = 8'b01100011;
DRAM[2200] = 8'b01100100;
DRAM[2201] = 8'b01101001;
DRAM[2202] = 8'b01101100;
DRAM[2203] = 8'b01101101;
DRAM[2204] = 8'b01110100;
DRAM[2205] = 8'b01110000;
DRAM[2206] = 8'b01110100;
DRAM[2207] = 8'b01110110;
DRAM[2208] = 8'b01110111;
DRAM[2209] = 8'b01111000;
DRAM[2210] = 8'b01111010;
DRAM[2211] = 8'b01111100;
DRAM[2212] = 8'b01111100;
DRAM[2213] = 8'b01111101;
DRAM[2214] = 8'b10000001;
DRAM[2215] = 8'b01110010;
DRAM[2216] = 8'b01110011;
DRAM[2217] = 8'b01111000;
DRAM[2218] = 8'b01110111;
DRAM[2219] = 8'b01110111;
DRAM[2220] = 8'b01111110;
DRAM[2221] = 8'b01111011;
DRAM[2222] = 8'b10000101;
DRAM[2223] = 8'b10000100;
DRAM[2224] = 8'b10000011;
DRAM[2225] = 8'b10001000;
DRAM[2226] = 8'b10000111;
DRAM[2227] = 8'b10000011;
DRAM[2228] = 8'b10001001;
DRAM[2229] = 8'b10001110;
DRAM[2230] = 8'b10010111;
DRAM[2231] = 8'b10100011;
DRAM[2232] = 8'b10101011;
DRAM[2233] = 8'b10101011;
DRAM[2234] = 8'b10110010;
DRAM[2235] = 8'b10110001;
DRAM[2236] = 8'b10110101;
DRAM[2237] = 8'b10110111;
DRAM[2238] = 8'b10111011;
DRAM[2239] = 8'b11000001;
DRAM[2240] = 8'b10111100;
DRAM[2241] = 8'b11000010;
DRAM[2242] = 8'b11000100;
DRAM[2243] = 8'b11000110;
DRAM[2244] = 8'b11000011;
DRAM[2245] = 8'b11001000;
DRAM[2246] = 8'b11000100;
DRAM[2247] = 8'b01111100;
DRAM[2248] = 8'b01100110;
DRAM[2249] = 8'b01101000;
DRAM[2250] = 8'b01101101;
DRAM[2251] = 8'b01110010;
DRAM[2252] = 8'b01110010;
DRAM[2253] = 8'b01101110;
DRAM[2254] = 8'b01101011;
DRAM[2255] = 8'b01101011;
DRAM[2256] = 8'b01101011;
DRAM[2257] = 8'b01100111;
DRAM[2258] = 8'b01101110;
DRAM[2259] = 8'b01111101;
DRAM[2260] = 8'b10001110;
DRAM[2261] = 8'b10011000;
DRAM[2262] = 8'b10010111;
DRAM[2263] = 8'b10011000;
DRAM[2264] = 8'b10010100;
DRAM[2265] = 8'b10001101;
DRAM[2266] = 8'b10001010;
DRAM[2267] = 8'b10001001;
DRAM[2268] = 8'b10001010;
DRAM[2269] = 8'b10010010;
DRAM[2270] = 8'b10010100;
DRAM[2271] = 8'b10001111;
DRAM[2272] = 8'b10001110;
DRAM[2273] = 8'b10010000;
DRAM[2274] = 8'b10010001;
DRAM[2275] = 8'b10001111;
DRAM[2276] = 8'b10001111;
DRAM[2277] = 8'b10001110;
DRAM[2278] = 8'b10001101;
DRAM[2279] = 8'b10010000;
DRAM[2280] = 8'b10001111;
DRAM[2281] = 8'b10010010;
DRAM[2282] = 8'b10010010;
DRAM[2283] = 8'b10010011;
DRAM[2284] = 8'b10010101;
DRAM[2285] = 8'b10011000;
DRAM[2286] = 8'b11000010;
DRAM[2287] = 8'b10001000;
DRAM[2288] = 8'b00101010;
DRAM[2289] = 8'b00101011;
DRAM[2290] = 8'b00101011;
DRAM[2291] = 8'b00101101;
DRAM[2292] = 8'b00101110;
DRAM[2293] = 8'b00110100;
DRAM[2294] = 8'b00110100;
DRAM[2295] = 8'b00110001;
DRAM[2296] = 8'b00110010;
DRAM[2297] = 8'b00110011;
DRAM[2298] = 8'b00110010;
DRAM[2299] = 8'b00101110;
DRAM[2300] = 8'b00110000;
DRAM[2301] = 8'b00111111;
DRAM[2302] = 8'b00101000;
DRAM[2303] = 8'b00100100;
DRAM[2304] = 8'b10101001;
DRAM[2305] = 8'b10100001;
DRAM[2306] = 8'b10001101;
DRAM[2307] = 8'b01101110;
DRAM[2308] = 8'b01001110;
DRAM[2309] = 8'b01010000;
DRAM[2310] = 8'b01101111;
DRAM[2311] = 8'b10001100;
DRAM[2312] = 8'b10011110;
DRAM[2313] = 8'b10101001;
DRAM[2314] = 8'b10100111;
DRAM[2315] = 8'b10100100;
DRAM[2316] = 8'b10100010;
DRAM[2317] = 8'b10011010;
DRAM[2318] = 8'b10001000;
DRAM[2319] = 8'b01101010;
DRAM[2320] = 8'b01001010;
DRAM[2321] = 8'b01001101;
DRAM[2322] = 8'b01011001;
DRAM[2323] = 8'b01100011;
DRAM[2324] = 8'b01100010;
DRAM[2325] = 8'b01100100;
DRAM[2326] = 8'b01100011;
DRAM[2327] = 8'b01100100;
DRAM[2328] = 8'b01100011;
DRAM[2329] = 8'b01100101;
DRAM[2330] = 8'b01101100;
DRAM[2331] = 8'b01101011;
DRAM[2332] = 8'b01101111;
DRAM[2333] = 8'b01110100;
DRAM[2334] = 8'b01110100;
DRAM[2335] = 8'b01110110;
DRAM[2336] = 8'b01111001;
DRAM[2337] = 8'b01110110;
DRAM[2338] = 8'b01111010;
DRAM[2339] = 8'b01111100;
DRAM[2340] = 8'b01111011;
DRAM[2341] = 8'b10000010;
DRAM[2342] = 8'b10010001;
DRAM[2343] = 8'b01110000;
DRAM[2344] = 8'b01110100;
DRAM[2345] = 8'b01101101;
DRAM[2346] = 8'b01110010;
DRAM[2347] = 8'b01110110;
DRAM[2348] = 8'b01111100;
DRAM[2349] = 8'b01111010;
DRAM[2350] = 8'b01111101;
DRAM[2351] = 8'b01111110;
DRAM[2352] = 8'b10000111;
DRAM[2353] = 8'b10001011;
DRAM[2354] = 8'b10000111;
DRAM[2355] = 8'b10000111;
DRAM[2356] = 8'b10001100;
DRAM[2357] = 8'b10001100;
DRAM[2358] = 8'b10010011;
DRAM[2359] = 8'b10011010;
DRAM[2360] = 8'b10100100;
DRAM[2361] = 8'b10101000;
DRAM[2362] = 8'b10101111;
DRAM[2363] = 8'b10110101;
DRAM[2364] = 8'b10110110;
DRAM[2365] = 8'b11000000;
DRAM[2366] = 8'b10111110;
DRAM[2367] = 8'b10111111;
DRAM[2368] = 8'b11000010;
DRAM[2369] = 8'b11000100;
DRAM[2370] = 8'b11000010;
DRAM[2371] = 8'b11000001;
DRAM[2372] = 8'b11000110;
DRAM[2373] = 8'b11000011;
DRAM[2374] = 8'b11000010;
DRAM[2375] = 8'b11001000;
DRAM[2376] = 8'b10001010;
DRAM[2377] = 8'b01101100;
DRAM[2378] = 8'b01011111;
DRAM[2379] = 8'b01101011;
DRAM[2380] = 8'b01101100;
DRAM[2381] = 8'b01101011;
DRAM[2382] = 8'b01101010;
DRAM[2383] = 8'b01101100;
DRAM[2384] = 8'b01101010;
DRAM[2385] = 8'b01100011;
DRAM[2386] = 8'b01101100;
DRAM[2387] = 8'b01111111;
DRAM[2388] = 8'b10010011;
DRAM[2389] = 8'b10011001;
DRAM[2390] = 8'b10011010;
DRAM[2391] = 8'b10011100;
DRAM[2392] = 8'b10010100;
DRAM[2393] = 8'b10001110;
DRAM[2394] = 8'b10000100;
DRAM[2395] = 8'b01111101;
DRAM[2396] = 8'b01111111;
DRAM[2397] = 8'b10001010;
DRAM[2398] = 8'b10010011;
DRAM[2399] = 8'b10010001;
DRAM[2400] = 8'b10001111;
DRAM[2401] = 8'b10010010;
DRAM[2402] = 8'b10010010;
DRAM[2403] = 8'b10010000;
DRAM[2404] = 8'b10001111;
DRAM[2405] = 8'b10001110;
DRAM[2406] = 8'b10001111;
DRAM[2407] = 8'b10010000;
DRAM[2408] = 8'b10010010;
DRAM[2409] = 8'b10010010;
DRAM[2410] = 8'b10010001;
DRAM[2411] = 8'b10010101;
DRAM[2412] = 8'b10010100;
DRAM[2413] = 8'b10011011;
DRAM[2414] = 8'b01110010;
DRAM[2415] = 8'b00101100;
DRAM[2416] = 8'b00101010;
DRAM[2417] = 8'b00101100;
DRAM[2418] = 8'b00110000;
DRAM[2419] = 8'b00110011;
DRAM[2420] = 8'b00110101;
DRAM[2421] = 8'b00110000;
DRAM[2422] = 8'b00101110;
DRAM[2423] = 8'b00101100;
DRAM[2424] = 8'b00110111;
DRAM[2425] = 8'b00110001;
DRAM[2426] = 8'b00101110;
DRAM[2427] = 8'b00110111;
DRAM[2428] = 8'b01000001;
DRAM[2429] = 8'b00110001;
DRAM[2430] = 8'b00100010;
DRAM[2431] = 8'b01110011;
DRAM[2432] = 8'b10100100;
DRAM[2433] = 8'b10010111;
DRAM[2434] = 8'b01111111;
DRAM[2435] = 8'b01011000;
DRAM[2436] = 8'b01011010;
DRAM[2437] = 8'b01010010;
DRAM[2438] = 8'b01110000;
DRAM[2439] = 8'b10001100;
DRAM[2440] = 8'b10011111;
DRAM[2441] = 8'b10100111;
DRAM[2442] = 8'b10101001;
DRAM[2443] = 8'b10100111;
DRAM[2444] = 8'b10100010;
DRAM[2445] = 8'b10011100;
DRAM[2446] = 8'b10001001;
DRAM[2447] = 8'b01101001;
DRAM[2448] = 8'b01001110;
DRAM[2449] = 8'b01010000;
DRAM[2450] = 8'b01011000;
DRAM[2451] = 8'b01100000;
DRAM[2452] = 8'b01100100;
DRAM[2453] = 8'b01100001;
DRAM[2454] = 8'b01100100;
DRAM[2455] = 8'b01100100;
DRAM[2456] = 8'b01100100;
DRAM[2457] = 8'b01100111;
DRAM[2458] = 8'b01101010;
DRAM[2459] = 8'b01101110;
DRAM[2460] = 8'b01110100;
DRAM[2461] = 8'b01110100;
DRAM[2462] = 8'b01110001;
DRAM[2463] = 8'b01110010;
DRAM[2464] = 8'b01110111;
DRAM[2465] = 8'b01111001;
DRAM[2466] = 8'b01111010;
DRAM[2467] = 8'b01111000;
DRAM[2468] = 8'b01111110;
DRAM[2469] = 8'b10001100;
DRAM[2470] = 8'b01110010;
DRAM[2471] = 8'b01101110;
DRAM[2472] = 8'b01101100;
DRAM[2473] = 8'b01110000;
DRAM[2474] = 8'b01111000;
DRAM[2475] = 8'b01110101;
DRAM[2476] = 8'b01111010;
DRAM[2477] = 8'b01111110;
DRAM[2478] = 8'b01111011;
DRAM[2479] = 8'b10000001;
DRAM[2480] = 8'b10000000;
DRAM[2481] = 8'b10000110;
DRAM[2482] = 8'b10000110;
DRAM[2483] = 8'b10000101;
DRAM[2484] = 8'b10001000;
DRAM[2485] = 8'b10010000;
DRAM[2486] = 8'b10001111;
DRAM[2487] = 8'b10010101;
DRAM[2488] = 8'b10100000;
DRAM[2489] = 8'b10101100;
DRAM[2490] = 8'b10110010;
DRAM[2491] = 8'b10111001;
DRAM[2492] = 8'b10111100;
DRAM[2493] = 8'b10111010;
DRAM[2494] = 8'b10111011;
DRAM[2495] = 8'b10111111;
DRAM[2496] = 8'b10111110;
DRAM[2497] = 8'b11000011;
DRAM[2498] = 8'b11000010;
DRAM[2499] = 8'b10111010;
DRAM[2500] = 8'b10111111;
DRAM[2501] = 8'b11000111;
DRAM[2502] = 8'b11010100;
DRAM[2503] = 8'b11011001;
DRAM[2504] = 8'b11100001;
DRAM[2505] = 8'b11100000;
DRAM[2506] = 8'b01110010;
DRAM[2507] = 8'b01011011;
DRAM[2508] = 8'b01101000;
DRAM[2509] = 8'b01100111;
DRAM[2510] = 8'b01100110;
DRAM[2511] = 8'b01101000;
DRAM[2512] = 8'b01100111;
DRAM[2513] = 8'b01100011;
DRAM[2514] = 8'b01101011;
DRAM[2515] = 8'b01111101;
DRAM[2516] = 8'b10001111;
DRAM[2517] = 8'b10011011;
DRAM[2518] = 8'b10011011;
DRAM[2519] = 8'b10011010;
DRAM[2520] = 8'b10010111;
DRAM[2521] = 8'b10010010;
DRAM[2522] = 8'b01111110;
DRAM[2523] = 8'b01101101;
DRAM[2524] = 8'b01101111;
DRAM[2525] = 8'b10000001;
DRAM[2526] = 8'b10001111;
DRAM[2527] = 8'b10010100;
DRAM[2528] = 8'b10010001;
DRAM[2529] = 8'b10010010;
DRAM[2530] = 8'b10010011;
DRAM[2531] = 8'b10001111;
DRAM[2532] = 8'b10001110;
DRAM[2533] = 8'b10001111;
DRAM[2534] = 8'b10001111;
DRAM[2535] = 8'b10010000;
DRAM[2536] = 8'b10001110;
DRAM[2537] = 8'b10010010;
DRAM[2538] = 8'b10010011;
DRAM[2539] = 8'b10010111;
DRAM[2540] = 8'b10011101;
DRAM[2541] = 8'b10000101;
DRAM[2542] = 8'b00111011;
DRAM[2543] = 8'b00101011;
DRAM[2544] = 8'b00101000;
DRAM[2545] = 8'b00101100;
DRAM[2546] = 8'b00110100;
DRAM[2547] = 8'b00110100;
DRAM[2548] = 8'b00110100;
DRAM[2549] = 8'b00101101;
DRAM[2550] = 8'b00101111;
DRAM[2551] = 8'b00110110;
DRAM[2552] = 8'b00110100;
DRAM[2553] = 8'b00101111;
DRAM[2554] = 8'b00110001;
DRAM[2555] = 8'b01000001;
DRAM[2556] = 8'b01000001;
DRAM[2557] = 8'b00100111;
DRAM[2558] = 8'b01011010;
DRAM[2559] = 8'b10100010;
DRAM[2560] = 8'b10011101;
DRAM[2561] = 8'b10001011;
DRAM[2562] = 8'b01101101;
DRAM[2563] = 8'b01010000;
DRAM[2564] = 8'b01010100;
DRAM[2565] = 8'b01010110;
DRAM[2566] = 8'b01110010;
DRAM[2567] = 8'b10001110;
DRAM[2568] = 8'b10011110;
DRAM[2569] = 8'b10100110;
DRAM[2570] = 8'b10100110;
DRAM[2571] = 8'b10100110;
DRAM[2572] = 8'b10100011;
DRAM[2573] = 8'b10011001;
DRAM[2574] = 8'b10000100;
DRAM[2575] = 8'b01100101;
DRAM[2576] = 8'b01001101;
DRAM[2577] = 8'b01001111;
DRAM[2578] = 8'b01011010;
DRAM[2579] = 8'b01011111;
DRAM[2580] = 8'b01100101;
DRAM[2581] = 8'b01100000;
DRAM[2582] = 8'b01100110;
DRAM[2583] = 8'b01100101;
DRAM[2584] = 8'b01100110;
DRAM[2585] = 8'b01101000;
DRAM[2586] = 8'b01101100;
DRAM[2587] = 8'b01101110;
DRAM[2588] = 8'b01110000;
DRAM[2589] = 8'b01110001;
DRAM[2590] = 8'b01110100;
DRAM[2591] = 8'b01110111;
DRAM[2592] = 8'b01111001;
DRAM[2593] = 8'b01111000;
DRAM[2594] = 8'b01111010;
DRAM[2595] = 8'b01111000;
DRAM[2596] = 8'b10000000;
DRAM[2597] = 8'b01111010;
DRAM[2598] = 8'b01101100;
DRAM[2599] = 8'b01110000;
DRAM[2600] = 8'b01110000;
DRAM[2601] = 8'b01110100;
DRAM[2602] = 8'b01110100;
DRAM[2603] = 8'b01111010;
DRAM[2604] = 8'b01111001;
DRAM[2605] = 8'b01110101;
DRAM[2606] = 8'b01111010;
DRAM[2607] = 8'b01111100;
DRAM[2608] = 8'b10000000;
DRAM[2609] = 8'b10000111;
DRAM[2610] = 8'b10000101;
DRAM[2611] = 8'b10000101;
DRAM[2612] = 8'b10000101;
DRAM[2613] = 8'b10001110;
DRAM[2614] = 8'b10001010;
DRAM[2615] = 8'b10010111;
DRAM[2616] = 8'b10011100;
DRAM[2617] = 8'b10101010;
DRAM[2618] = 8'b10110111;
DRAM[2619] = 8'b10111001;
DRAM[2620] = 8'b10111011;
DRAM[2621] = 8'b10111010;
DRAM[2622] = 8'b10111011;
DRAM[2623] = 8'b10111101;
DRAM[2624] = 8'b10111001;
DRAM[2625] = 8'b10110101;
DRAM[2626] = 8'b11000001;
DRAM[2627] = 8'b11010001;
DRAM[2628] = 8'b11010100;
DRAM[2629] = 8'b11010010;
DRAM[2630] = 8'b11010100;
DRAM[2631] = 8'b11010011;
DRAM[2632] = 8'b11011000;
DRAM[2633] = 8'b11100001;
DRAM[2634] = 8'b11000110;
DRAM[2635] = 8'b01010011;
DRAM[2636] = 8'b01011011;
DRAM[2637] = 8'b01100101;
DRAM[2638] = 8'b01100100;
DRAM[2639] = 8'b01100101;
DRAM[2640] = 8'b01100011;
DRAM[2641] = 8'b01011101;
DRAM[2642] = 8'b01101010;
DRAM[2643] = 8'b01111010;
DRAM[2644] = 8'b10001111;
DRAM[2645] = 8'b10011000;
DRAM[2646] = 8'b10011010;
DRAM[2647] = 8'b10011010;
DRAM[2648] = 8'b10011011;
DRAM[2649] = 8'b10010011;
DRAM[2650] = 8'b10000001;
DRAM[2651] = 8'b01100000;
DRAM[2652] = 8'b01010100;
DRAM[2653] = 8'b01101100;
DRAM[2654] = 8'b10000111;
DRAM[2655] = 8'b10010001;
DRAM[2656] = 8'b10010001;
DRAM[2657] = 8'b10001111;
DRAM[2658] = 8'b10010011;
DRAM[2659] = 8'b10001111;
DRAM[2660] = 8'b10001110;
DRAM[2661] = 8'b10001111;
DRAM[2662] = 8'b10001110;
DRAM[2663] = 8'b10010011;
DRAM[2664] = 8'b10010011;
DRAM[2665] = 8'b10010010;
DRAM[2666] = 8'b10010101;
DRAM[2667] = 8'b10011000;
DRAM[2668] = 8'b10010100;
DRAM[2669] = 8'b01000011;
DRAM[2670] = 8'b00101100;
DRAM[2671] = 8'b00100111;
DRAM[2672] = 8'b00101110;
DRAM[2673] = 8'b00110011;
DRAM[2674] = 8'b00110111;
DRAM[2675] = 8'b00110100;
DRAM[2676] = 8'b00101111;
DRAM[2677] = 8'b00101010;
DRAM[2678] = 8'b00110110;
DRAM[2679] = 8'b00110100;
DRAM[2680] = 8'b00101101;
DRAM[2681] = 8'b00101110;
DRAM[2682] = 8'b00111010;
DRAM[2683] = 8'b01001101;
DRAM[2684] = 8'b00110111;
DRAM[2685] = 8'b01010110;
DRAM[2686] = 8'b10010001;
DRAM[2687] = 8'b10100010;
DRAM[2688] = 8'b10010100;
DRAM[2689] = 8'b01111001;
DRAM[2690] = 8'b01010100;
DRAM[2691] = 8'b01011000;
DRAM[2692] = 8'b01010110;
DRAM[2693] = 8'b01011000;
DRAM[2694] = 8'b01110010;
DRAM[2695] = 8'b10001011;
DRAM[2696] = 8'b10011110;
DRAM[2697] = 8'b10100111;
DRAM[2698] = 8'b10101000;
DRAM[2699] = 8'b10100101;
DRAM[2700] = 8'b10100011;
DRAM[2701] = 8'b10011001;
DRAM[2702] = 8'b10000101;
DRAM[2703] = 8'b01101011;
DRAM[2704] = 8'b01010000;
DRAM[2705] = 8'b01010010;
DRAM[2706] = 8'b01011001;
DRAM[2707] = 8'b01011110;
DRAM[2708] = 8'b01100010;
DRAM[2709] = 8'b01100010;
DRAM[2710] = 8'b01100101;
DRAM[2711] = 8'b01101001;
DRAM[2712] = 8'b01100100;
DRAM[2713] = 8'b01100110;
DRAM[2714] = 8'b01101011;
DRAM[2715] = 8'b01110000;
DRAM[2716] = 8'b01110010;
DRAM[2717] = 8'b01110010;
DRAM[2718] = 8'b01110101;
DRAM[2719] = 8'b01111000;
DRAM[2720] = 8'b01111000;
DRAM[2721] = 8'b01111001;
DRAM[2722] = 8'b01111100;
DRAM[2723] = 8'b01111100;
DRAM[2724] = 8'b01111011;
DRAM[2725] = 8'b01101011;
DRAM[2726] = 8'b01101110;
DRAM[2727] = 8'b01110000;
DRAM[2728] = 8'b01110100;
DRAM[2729] = 8'b01110101;
DRAM[2730] = 8'b01111100;
DRAM[2731] = 8'b01111001;
DRAM[2732] = 8'b01110111;
DRAM[2733] = 8'b01110111;
DRAM[2734] = 8'b01111001;
DRAM[2735] = 8'b10000010;
DRAM[2736] = 8'b10000001;
DRAM[2737] = 8'b10001101;
DRAM[2738] = 8'b10001001;
DRAM[2739] = 8'b10001001;
DRAM[2740] = 8'b10000111;
DRAM[2741] = 8'b10001111;
DRAM[2742] = 8'b10001110;
DRAM[2743] = 8'b10010111;
DRAM[2744] = 8'b10011111;
DRAM[2745] = 8'b10101001;
DRAM[2746] = 8'b10110100;
DRAM[2747] = 8'b10110111;
DRAM[2748] = 8'b10111001;
DRAM[2749] = 8'b10111101;
DRAM[2750] = 8'b10101111;
DRAM[2751] = 8'b10101110;
DRAM[2752] = 8'b11000000;
DRAM[2753] = 8'b11010001;
DRAM[2754] = 8'b11010010;
DRAM[2755] = 8'b11001110;
DRAM[2756] = 8'b11010000;
DRAM[2757] = 8'b11001111;
DRAM[2758] = 8'b11010000;
DRAM[2759] = 8'b11010011;
DRAM[2760] = 8'b11010010;
DRAM[2761] = 8'b11011010;
DRAM[2762] = 8'b11011110;
DRAM[2763] = 8'b10100101;
DRAM[2764] = 8'b01001110;
DRAM[2765] = 8'b01011001;
DRAM[2766] = 8'b01100000;
DRAM[2767] = 8'b01100011;
DRAM[2768] = 8'b01100010;
DRAM[2769] = 8'b01011111;
DRAM[2770] = 8'b01100111;
DRAM[2771] = 8'b01111010;
DRAM[2772] = 8'b10001101;
DRAM[2773] = 8'b10011000;
DRAM[2774] = 8'b10011001;
DRAM[2775] = 8'b10011000;
DRAM[2776] = 8'b10011010;
DRAM[2777] = 8'b10010010;
DRAM[2778] = 8'b10000101;
DRAM[2779] = 8'b01011110;
DRAM[2780] = 8'b00111001;
DRAM[2781] = 8'b01010000;
DRAM[2782] = 8'b01111010;
DRAM[2783] = 8'b10001011;
DRAM[2784] = 8'b10010101;
DRAM[2785] = 8'b10010010;
DRAM[2786] = 8'b10010010;
DRAM[2787] = 8'b10010001;
DRAM[2788] = 8'b10001111;
DRAM[2789] = 8'b10001110;
DRAM[2790] = 8'b10001111;
DRAM[2791] = 8'b10010000;
DRAM[2792] = 8'b10001110;
DRAM[2793] = 8'b10010010;
DRAM[2794] = 8'b10010111;
DRAM[2795] = 8'b10011010;
DRAM[2796] = 8'b01100010;
DRAM[2797] = 8'b00101001;
DRAM[2798] = 8'b00101001;
DRAM[2799] = 8'b00101010;
DRAM[2800] = 8'b00110100;
DRAM[2801] = 8'b00110100;
DRAM[2802] = 8'b00110100;
DRAM[2803] = 8'b00110110;
DRAM[2804] = 8'b00101010;
DRAM[2805] = 8'b00110011;
DRAM[2806] = 8'b00110100;
DRAM[2807] = 8'b00101101;
DRAM[2808] = 8'b00110000;
DRAM[2809] = 8'b00111111;
DRAM[2810] = 8'b01001000;
DRAM[2811] = 8'b01000101;
DRAM[2812] = 8'b01011010;
DRAM[2813] = 8'b10001010;
DRAM[2814] = 8'b10010100;
DRAM[2815] = 8'b10010111;
DRAM[2816] = 8'b10000100;
DRAM[2817] = 8'b01100000;
DRAM[2818] = 8'b01010100;
DRAM[2819] = 8'b01011000;
DRAM[2820] = 8'b01010110;
DRAM[2821] = 8'b01011000;
DRAM[2822] = 8'b01110000;
DRAM[2823] = 8'b10001110;
DRAM[2824] = 8'b10011011;
DRAM[2825] = 8'b10100101;
DRAM[2826] = 8'b10100111;
DRAM[2827] = 8'b10100110;
DRAM[2828] = 8'b10100010;
DRAM[2829] = 8'b10011000;
DRAM[2830] = 8'b10000111;
DRAM[2831] = 8'b01101000;
DRAM[2832] = 8'b01001101;
DRAM[2833] = 8'b01010010;
DRAM[2834] = 8'b01011011;
DRAM[2835] = 8'b01100010;
DRAM[2836] = 8'b01100010;
DRAM[2837] = 8'b01100101;
DRAM[2838] = 8'b01100011;
DRAM[2839] = 8'b01100101;
DRAM[2840] = 8'b01100100;
DRAM[2841] = 8'b01100101;
DRAM[2842] = 8'b01101100;
DRAM[2843] = 8'b01101100;
DRAM[2844] = 8'b01110100;
DRAM[2845] = 8'b01110101;
DRAM[2846] = 8'b01110101;
DRAM[2847] = 8'b01110111;
DRAM[2848] = 8'b01111001;
DRAM[2849] = 8'b01111001;
DRAM[2850] = 8'b01111011;
DRAM[2851] = 8'b01111110;
DRAM[2852] = 8'b01101101;
DRAM[2853] = 8'b01101001;
DRAM[2854] = 8'b01101111;
DRAM[2855] = 8'b01110010;
DRAM[2856] = 8'b01110010;
DRAM[2857] = 8'b01110101;
DRAM[2858] = 8'b01110110;
DRAM[2859] = 8'b01110111;
DRAM[2860] = 8'b01110001;
DRAM[2861] = 8'b01111001;
DRAM[2862] = 8'b01111101;
DRAM[2863] = 8'b01111110;
DRAM[2864] = 8'b10001001;
DRAM[2865] = 8'b10000110;
DRAM[2866] = 8'b10001000;
DRAM[2867] = 8'b10001011;
DRAM[2868] = 8'b10001110;
DRAM[2869] = 8'b10001110;
DRAM[2870] = 8'b10010101;
DRAM[2871] = 8'b10010000;
DRAM[2872] = 8'b10011101;
DRAM[2873] = 8'b10100000;
DRAM[2874] = 8'b10110010;
DRAM[2875] = 8'b10110001;
DRAM[2876] = 8'b10110110;
DRAM[2877] = 8'b10100001;
DRAM[2878] = 8'b10111010;
DRAM[2879] = 8'b11001100;
DRAM[2880] = 8'b11010010;
DRAM[2881] = 8'b11001101;
DRAM[2882] = 8'b11001110;
DRAM[2883] = 8'b11001100;
DRAM[2884] = 8'b11010000;
DRAM[2885] = 8'b11001111;
DRAM[2886] = 8'b11001100;
DRAM[2887] = 8'b11001100;
DRAM[2888] = 8'b11010001;
DRAM[2889] = 8'b11010011;
DRAM[2890] = 8'b11011110;
DRAM[2891] = 8'b11011110;
DRAM[2892] = 8'b10000100;
DRAM[2893] = 8'b01001110;
DRAM[2894] = 8'b01010111;
DRAM[2895] = 8'b01011100;
DRAM[2896] = 8'b01011110;
DRAM[2897] = 8'b01011110;
DRAM[2898] = 8'b01100110;
DRAM[2899] = 8'b01111010;
DRAM[2900] = 8'b10001100;
DRAM[2901] = 8'b10011001;
DRAM[2902] = 8'b10011100;
DRAM[2903] = 8'b10011010;
DRAM[2904] = 8'b10011000;
DRAM[2905] = 8'b10010110;
DRAM[2906] = 8'b10000110;
DRAM[2907] = 8'b01100010;
DRAM[2908] = 8'b00110100;
DRAM[2909] = 8'b00111010;
DRAM[2910] = 8'b01100101;
DRAM[2911] = 8'b10000001;
DRAM[2912] = 8'b10010001;
DRAM[2913] = 8'b10010101;
DRAM[2914] = 8'b10010001;
DRAM[2915] = 8'b10010000;
DRAM[2916] = 8'b10001110;
DRAM[2917] = 8'b10001111;
DRAM[2918] = 8'b10010001;
DRAM[2919] = 8'b10010010;
DRAM[2920] = 8'b10010001;
DRAM[2921] = 8'b10010100;
DRAM[2922] = 8'b10011001;
DRAM[2923] = 8'b01111011;
DRAM[2924] = 8'b00110001;
DRAM[2925] = 8'b00111000;
DRAM[2926] = 8'b00101110;
DRAM[2927] = 8'b00110011;
DRAM[2928] = 8'b00110110;
DRAM[2929] = 8'b00110111;
DRAM[2930] = 8'b00110100;
DRAM[2931] = 8'b00101110;
DRAM[2932] = 8'b00110001;
DRAM[2933] = 8'b00111010;
DRAM[2934] = 8'b00101110;
DRAM[2935] = 8'b00110011;
DRAM[2936] = 8'b00111010;
DRAM[2937] = 8'b01000010;
DRAM[2938] = 8'b01001000;
DRAM[2939] = 8'b01011011;
DRAM[2940] = 8'b10000101;
DRAM[2941] = 8'b10010111;
DRAM[2942] = 8'b10001110;
DRAM[2943] = 8'b10001111;
DRAM[2944] = 8'b01101110;
DRAM[2945] = 8'b01010110;
DRAM[2946] = 8'b01011000;
DRAM[2947] = 8'b01011010;
DRAM[2948] = 8'b01011000;
DRAM[2949] = 8'b01010111;
DRAM[2950] = 8'b01101111;
DRAM[2951] = 8'b10001101;
DRAM[2952] = 8'b10011100;
DRAM[2953] = 8'b10100011;
DRAM[2954] = 8'b10101001;
DRAM[2955] = 8'b10100101;
DRAM[2956] = 8'b10100011;
DRAM[2957] = 8'b10011010;
DRAM[2958] = 8'b10000100;
DRAM[2959] = 8'b01101000;
DRAM[2960] = 8'b01001101;
DRAM[2961] = 8'b01010010;
DRAM[2962] = 8'b01011100;
DRAM[2963] = 8'b01100000;
DRAM[2964] = 8'b01100000;
DRAM[2965] = 8'b01100010;
DRAM[2966] = 8'b01100011;
DRAM[2967] = 8'b01100101;
DRAM[2968] = 8'b01100100;
DRAM[2969] = 8'b01101001;
DRAM[2970] = 8'b01101000;
DRAM[2971] = 8'b01101111;
DRAM[2972] = 8'b01110011;
DRAM[2973] = 8'b01110110;
DRAM[2974] = 8'b01110100;
DRAM[2975] = 8'b01110111;
DRAM[2976] = 8'b01110111;
DRAM[2977] = 8'b01111011;
DRAM[2978] = 8'b01111101;
DRAM[2979] = 8'b01110010;
DRAM[2980] = 8'b01101011;
DRAM[2981] = 8'b01110000;
DRAM[2982] = 8'b01110010;
DRAM[2983] = 8'b01110010;
DRAM[2984] = 8'b01110110;
DRAM[2985] = 8'b01110111;
DRAM[2986] = 8'b01110000;
DRAM[2987] = 8'b01101110;
DRAM[2988] = 8'b01110110;
DRAM[2989] = 8'b01111101;
DRAM[2990] = 8'b10000010;
DRAM[2991] = 8'b10000001;
DRAM[2992] = 8'b10001011;
DRAM[2993] = 8'b10001011;
DRAM[2994] = 8'b10010000;
DRAM[2995] = 8'b10010001;
DRAM[2996] = 8'b10010010;
DRAM[2997] = 8'b10001010;
DRAM[2998] = 8'b10001010;
DRAM[2999] = 8'b10010011;
DRAM[3000] = 8'b10011011;
DRAM[3001] = 8'b10101000;
DRAM[3002] = 8'b10100110;
DRAM[3003] = 8'b10011100;
DRAM[3004] = 8'b10101000;
DRAM[3005] = 8'b11001101;
DRAM[3006] = 8'b11001110;
DRAM[3007] = 8'b11001000;
DRAM[3008] = 8'b11001010;
DRAM[3009] = 8'b11010011;
DRAM[3010] = 8'b11001110;
DRAM[3011] = 8'b11001000;
DRAM[3012] = 8'b11000011;
DRAM[3013] = 8'b11001001;
DRAM[3014] = 8'b11001011;
DRAM[3015] = 8'b11010100;
DRAM[3016] = 8'b11010011;
DRAM[3017] = 8'b11010010;
DRAM[3018] = 8'b11010111;
DRAM[3019] = 8'b11011110;
DRAM[3020] = 8'b11011001;
DRAM[3021] = 8'b01010100;
DRAM[3022] = 8'b01001100;
DRAM[3023] = 8'b01010010;
DRAM[3024] = 8'b01011000;
DRAM[3025] = 8'b01011010;
DRAM[3026] = 8'b01100100;
DRAM[3027] = 8'b01111011;
DRAM[3028] = 8'b10001110;
DRAM[3029] = 8'b10011001;
DRAM[3030] = 8'b10011010;
DRAM[3031] = 8'b10011001;
DRAM[3032] = 8'b10011010;
DRAM[3033] = 8'b10010101;
DRAM[3034] = 8'b10001001;
DRAM[3035] = 8'b01100111;
DRAM[3036] = 8'b00110000;
DRAM[3037] = 8'b00110000;
DRAM[3038] = 8'b01010111;
DRAM[3039] = 8'b01110001;
DRAM[3040] = 8'b10001010;
DRAM[3041] = 8'b10010010;
DRAM[3042] = 8'b10010010;
DRAM[3043] = 8'b10010001;
DRAM[3044] = 8'b10001110;
DRAM[3045] = 8'b10001101;
DRAM[3046] = 8'b10010000;
DRAM[3047] = 8'b10010010;
DRAM[3048] = 8'b10010010;
DRAM[3049] = 8'b10010111;
DRAM[3050] = 8'b10010101;
DRAM[3051] = 8'b00111011;
DRAM[3052] = 8'b00101010;
DRAM[3053] = 8'b00101010;
DRAM[3054] = 8'b00110000;
DRAM[3055] = 8'b00110110;
DRAM[3056] = 8'b00110100;
DRAM[3057] = 8'b00110100;
DRAM[3058] = 8'b00101011;
DRAM[3059] = 8'b00101110;
DRAM[3060] = 8'b00111010;
DRAM[3061] = 8'b00110011;
DRAM[3062] = 8'b00110100;
DRAM[3063] = 8'b00110001;
DRAM[3064] = 8'b00110111;
DRAM[3065] = 8'b01000101;
DRAM[3066] = 8'b01011100;
DRAM[3067] = 8'b10000010;
DRAM[3068] = 8'b10010011;
DRAM[3069] = 8'b10010100;
DRAM[3070] = 8'b10001110;
DRAM[3071] = 8'b10100010;
DRAM[3072] = 8'b01011000;
DRAM[3073] = 8'b01010110;
DRAM[3074] = 8'b01011011;
DRAM[3075] = 8'b01011100;
DRAM[3076] = 8'b01011011;
DRAM[3077] = 8'b01010110;
DRAM[3078] = 8'b01110000;
DRAM[3079] = 8'b10001000;
DRAM[3080] = 8'b10011010;
DRAM[3081] = 8'b10100011;
DRAM[3082] = 8'b10100111;
DRAM[3083] = 8'b10100100;
DRAM[3084] = 8'b10100010;
DRAM[3085] = 8'b10011011;
DRAM[3086] = 8'b10000101;
DRAM[3087] = 8'b01100111;
DRAM[3088] = 8'b01001101;
DRAM[3089] = 8'b01001110;
DRAM[3090] = 8'b01011101;
DRAM[3091] = 8'b01100000;
DRAM[3092] = 8'b01100010;
DRAM[3093] = 8'b01100101;
DRAM[3094] = 8'b01100000;
DRAM[3095] = 8'b01100011;
DRAM[3096] = 8'b01100100;
DRAM[3097] = 8'b01100110;
DRAM[3098] = 8'b01101001;
DRAM[3099] = 8'b01101100;
DRAM[3100] = 8'b01110010;
DRAM[3101] = 8'b01110100;
DRAM[3102] = 8'b01110010;
DRAM[3103] = 8'b01110110;
DRAM[3104] = 8'b01111001;
DRAM[3105] = 8'b01111110;
DRAM[3106] = 8'b01110111;
DRAM[3107] = 8'b01110010;
DRAM[3108] = 8'b01110100;
DRAM[3109] = 8'b01101110;
DRAM[3110] = 8'b01101110;
DRAM[3111] = 8'b01110101;
DRAM[3112] = 8'b01110111;
DRAM[3113] = 8'b01110001;
DRAM[3114] = 8'b01110110;
DRAM[3115] = 8'b01111000;
DRAM[3116] = 8'b01110111;
DRAM[3117] = 8'b10000000;
DRAM[3118] = 8'b01111110;
DRAM[3119] = 8'b10000110;
DRAM[3120] = 8'b10001010;
DRAM[3121] = 8'b10001010;
DRAM[3122] = 8'b10001100;
DRAM[3123] = 8'b10001111;
DRAM[3124] = 8'b10001001;
DRAM[3125] = 8'b10001100;
DRAM[3126] = 8'b10001100;
DRAM[3127] = 8'b10010000;
DRAM[3128] = 8'b10011111;
DRAM[3129] = 8'b10100100;
DRAM[3130] = 8'b10001111;
DRAM[3131] = 8'b10110101;
DRAM[3132] = 8'b11000100;
DRAM[3133] = 8'b11001001;
DRAM[3134] = 8'b11001001;
DRAM[3135] = 8'b11001110;
DRAM[3136] = 8'b11001000;
DRAM[3137] = 8'b11001001;
DRAM[3138] = 8'b11000011;
DRAM[3139] = 8'b11000100;
DRAM[3140] = 8'b11001101;
DRAM[3141] = 8'b11001001;
DRAM[3142] = 8'b11001000;
DRAM[3143] = 8'b11001001;
DRAM[3144] = 8'b11001100;
DRAM[3145] = 8'b11010001;
DRAM[3146] = 8'b11010100;
DRAM[3147] = 8'b11010101;
DRAM[3148] = 8'b11011010;
DRAM[3149] = 8'b11010111;
DRAM[3150] = 8'b10010000;
DRAM[3151] = 8'b01001010;
DRAM[3152] = 8'b01001110;
DRAM[3153] = 8'b01010110;
DRAM[3154] = 8'b01100100;
DRAM[3155] = 8'b01111100;
DRAM[3156] = 8'b10001111;
DRAM[3157] = 8'b10011000;
DRAM[3158] = 8'b10011011;
DRAM[3159] = 8'b10011011;
DRAM[3160] = 8'b10011001;
DRAM[3161] = 8'b10011000;
DRAM[3162] = 8'b10001000;
DRAM[3163] = 8'b01100100;
DRAM[3164] = 8'b00110100;
DRAM[3165] = 8'b00101100;
DRAM[3166] = 8'b00111101;
DRAM[3167] = 8'b01100010;
DRAM[3168] = 8'b01111110;
DRAM[3169] = 8'b10001110;
DRAM[3170] = 8'b10010110;
DRAM[3171] = 8'b10010000;
DRAM[3172] = 8'b10001111;
DRAM[3173] = 8'b10001110;
DRAM[3174] = 8'b10010001;
DRAM[3175] = 8'b10010001;
DRAM[3176] = 8'b10010111;
DRAM[3177] = 8'b10011001;
DRAM[3178] = 8'b01100011;
DRAM[3179] = 8'b00101001;
DRAM[3180] = 8'b00100110;
DRAM[3181] = 8'b00101010;
DRAM[3182] = 8'b00111000;
DRAM[3183] = 8'b00111001;
DRAM[3184] = 8'b00110011;
DRAM[3185] = 8'b00101110;
DRAM[3186] = 8'b00101010;
DRAM[3187] = 8'b00111000;
DRAM[3188] = 8'b00110001;
DRAM[3189] = 8'b00101110;
DRAM[3190] = 8'b00110100;
DRAM[3191] = 8'b00110110;
DRAM[3192] = 8'b01000001;
DRAM[3193] = 8'b01001101;
DRAM[3194] = 8'b01111111;
DRAM[3195] = 8'b10010001;
DRAM[3196] = 8'b10010101;
DRAM[3197] = 8'b10001101;
DRAM[3198] = 8'b10100000;
DRAM[3199] = 8'b10100101;
DRAM[3200] = 8'b01011000;
DRAM[3201] = 8'b01011100;
DRAM[3202] = 8'b01011010;
DRAM[3203] = 8'b01011010;
DRAM[3204] = 8'b01011000;
DRAM[3205] = 8'b01011010;
DRAM[3206] = 8'b01101100;
DRAM[3207] = 8'b10001011;
DRAM[3208] = 8'b10011010;
DRAM[3209] = 8'b10100100;
DRAM[3210] = 8'b10100101;
DRAM[3211] = 8'b10100110;
DRAM[3212] = 8'b10100010;
DRAM[3213] = 8'b10011001;
DRAM[3214] = 8'b10000101;
DRAM[3215] = 8'b01101001;
DRAM[3216] = 8'b01001110;
DRAM[3217] = 8'b01001110;
DRAM[3218] = 8'b01011000;
DRAM[3219] = 8'b01011110;
DRAM[3220] = 8'b01100100;
DRAM[3221] = 8'b01100010;
DRAM[3222] = 8'b01100110;
DRAM[3223] = 8'b01100100;
DRAM[3224] = 8'b01101000;
DRAM[3225] = 8'b01100100;
DRAM[3226] = 8'b01101010;
DRAM[3227] = 8'b01101111;
DRAM[3228] = 8'b01110010;
DRAM[3229] = 8'b01110011;
DRAM[3230] = 8'b01111000;
DRAM[3231] = 8'b01110101;
DRAM[3232] = 8'b01110110;
DRAM[3233] = 8'b10000010;
DRAM[3234] = 8'b01101110;
DRAM[3235] = 8'b01101000;
DRAM[3236] = 8'b01110010;
DRAM[3237] = 8'b01110011;
DRAM[3238] = 8'b01110001;
DRAM[3239] = 8'b01110001;
DRAM[3240] = 8'b01101111;
DRAM[3241] = 8'b01110011;
DRAM[3242] = 8'b01110100;
DRAM[3243] = 8'b01111001;
DRAM[3244] = 8'b10000101;
DRAM[3245] = 8'b01111110;
DRAM[3246] = 8'b10000110;
DRAM[3247] = 8'b10001010;
DRAM[3248] = 8'b10001101;
DRAM[3249] = 8'b10001001;
DRAM[3250] = 8'b10001011;
DRAM[3251] = 8'b10001101;
DRAM[3252] = 8'b10000101;
DRAM[3253] = 8'b10000110;
DRAM[3254] = 8'b10001110;
DRAM[3255] = 8'b10001001;
DRAM[3256] = 8'b10001110;
DRAM[3257] = 8'b10010110;
DRAM[3258] = 8'b10111111;
DRAM[3259] = 8'b11000101;
DRAM[3260] = 8'b11000100;
DRAM[3261] = 8'b11000100;
DRAM[3262] = 8'b11000100;
DRAM[3263] = 8'b11000100;
DRAM[3264] = 8'b11000101;
DRAM[3265] = 8'b11000111;
DRAM[3266] = 8'b11000110;
DRAM[3267] = 8'b11000101;
DRAM[3268] = 8'b11001000;
DRAM[3269] = 8'b11001110;
DRAM[3270] = 8'b11001110;
DRAM[3271] = 8'b11001111;
DRAM[3272] = 8'b11001111;
DRAM[3273] = 8'b11001111;
DRAM[3274] = 8'b11010001;
DRAM[3275] = 8'b11010000;
DRAM[3276] = 8'b11010110;
DRAM[3277] = 8'b11010111;
DRAM[3278] = 8'b11011111;
DRAM[3279] = 8'b10001101;
DRAM[3280] = 8'b01000010;
DRAM[3281] = 8'b01001011;
DRAM[3282] = 8'b01011110;
DRAM[3283] = 8'b01111010;
DRAM[3284] = 8'b10001101;
DRAM[3285] = 8'b10011010;
DRAM[3286] = 8'b10011001;
DRAM[3287] = 8'b10011010;
DRAM[3288] = 8'b10011000;
DRAM[3289] = 8'b10010111;
DRAM[3290] = 8'b10000110;
DRAM[3291] = 8'b01100110;
DRAM[3292] = 8'b00111011;
DRAM[3293] = 8'b00101101;
DRAM[3294] = 8'b00101110;
DRAM[3295] = 8'b01000101;
DRAM[3296] = 8'b01101100;
DRAM[3297] = 8'b10000110;
DRAM[3298] = 8'b10010011;
DRAM[3299] = 8'b10010001;
DRAM[3300] = 8'b10001100;
DRAM[3301] = 8'b10001101;
DRAM[3302] = 8'b10010000;
DRAM[3303] = 8'b10010011;
DRAM[3304] = 8'b10011000;
DRAM[3305] = 8'b10000000;
DRAM[3306] = 8'b00101101;
DRAM[3307] = 8'b00101010;
DRAM[3308] = 8'b00101010;
DRAM[3309] = 8'b00101111;
DRAM[3310] = 8'b00110110;
DRAM[3311] = 8'b00110111;
DRAM[3312] = 8'b00110110;
DRAM[3313] = 8'b00101110;
DRAM[3314] = 8'b00110001;
DRAM[3315] = 8'b00110100;
DRAM[3316] = 8'b00101111;
DRAM[3317] = 8'b00110010;
DRAM[3318] = 8'b00110100;
DRAM[3319] = 8'b00111000;
DRAM[3320] = 8'b01000001;
DRAM[3321] = 8'b01111000;
DRAM[3322] = 8'b10001111;
DRAM[3323] = 8'b10010001;
DRAM[3324] = 8'b10010000;
DRAM[3325] = 8'b10011111;
DRAM[3326] = 8'b10100100;
DRAM[3327] = 8'b10100100;
DRAM[3328] = 8'b01010101;
DRAM[3329] = 8'b01100000;
DRAM[3330] = 8'b01011100;
DRAM[3331] = 8'b01011100;
DRAM[3332] = 8'b01011011;
DRAM[3333] = 8'b01011010;
DRAM[3334] = 8'b01110000;
DRAM[3335] = 8'b10001001;
DRAM[3336] = 8'b10011000;
DRAM[3337] = 8'b10100011;
DRAM[3338] = 8'b10100011;
DRAM[3339] = 8'b10100001;
DRAM[3340] = 8'b10100000;
DRAM[3341] = 8'b10011001;
DRAM[3342] = 8'b10000111;
DRAM[3343] = 8'b01100110;
DRAM[3344] = 8'b01010010;
DRAM[3345] = 8'b01001110;
DRAM[3346] = 8'b01011010;
DRAM[3347] = 8'b01011100;
DRAM[3348] = 8'b01011111;
DRAM[3349] = 8'b01100010;
DRAM[3350] = 8'b01100111;
DRAM[3351] = 8'b01100010;
DRAM[3352] = 8'b01100100;
DRAM[3353] = 8'b01100101;
DRAM[3354] = 8'b01101000;
DRAM[3355] = 8'b01101110;
DRAM[3356] = 8'b01110000;
DRAM[3357] = 8'b01110101;
DRAM[3358] = 8'b01110101;
DRAM[3359] = 8'b01101111;
DRAM[3360] = 8'b10001101;
DRAM[3361] = 8'b10000000;
DRAM[3362] = 8'b01101000;
DRAM[3363] = 8'b01101000;
DRAM[3364] = 8'b01101100;
DRAM[3365] = 8'b01110001;
DRAM[3366] = 8'b01110001;
DRAM[3367] = 8'b01110001;
DRAM[3368] = 8'b01110011;
DRAM[3369] = 8'b01110000;
DRAM[3370] = 8'b01111001;
DRAM[3371] = 8'b01111001;
DRAM[3372] = 8'b10000101;
DRAM[3373] = 8'b10001000;
DRAM[3374] = 8'b10010000;
DRAM[3375] = 8'b10001100;
DRAM[3376] = 8'b10000111;
DRAM[3377] = 8'b10001101;
DRAM[3378] = 8'b10001100;
DRAM[3379] = 8'b10001001;
DRAM[3380] = 8'b10000011;
DRAM[3381] = 8'b10000000;
DRAM[3382] = 8'b10000101;
DRAM[3383] = 8'b10000100;
DRAM[3384] = 8'b10101100;
DRAM[3385] = 8'b10110010;
DRAM[3386] = 8'b11000010;
DRAM[3387] = 8'b11000111;
DRAM[3388] = 8'b11000000;
DRAM[3389] = 8'b11000001;
DRAM[3390] = 8'b10111110;
DRAM[3391] = 8'b10111101;
DRAM[3392] = 8'b10111111;
DRAM[3393] = 8'b11000101;
DRAM[3394] = 8'b11001110;
DRAM[3395] = 8'b11001010;
DRAM[3396] = 8'b11001101;
DRAM[3397] = 8'b11001011;
DRAM[3398] = 8'b11001111;
DRAM[3399] = 8'b11001101;
DRAM[3400] = 8'b11010000;
DRAM[3401] = 8'b11001111;
DRAM[3402] = 8'b11010001;
DRAM[3403] = 8'b11001111;
DRAM[3404] = 8'b11010011;
DRAM[3405] = 8'b11010110;
DRAM[3406] = 8'b11011000;
DRAM[3407] = 8'b11011101;
DRAM[3408] = 8'b01100001;
DRAM[3409] = 8'b01000100;
DRAM[3410] = 8'b01011000;
DRAM[3411] = 8'b01110111;
DRAM[3412] = 8'b10001011;
DRAM[3413] = 8'b10010111;
DRAM[3414] = 8'b10011001;
DRAM[3415] = 8'b10011010;
DRAM[3416] = 8'b10011001;
DRAM[3417] = 8'b10011000;
DRAM[3418] = 8'b10000111;
DRAM[3419] = 8'b01101010;
DRAM[3420] = 8'b00111000;
DRAM[3421] = 8'b00101100;
DRAM[3422] = 8'b00101101;
DRAM[3423] = 8'b00101110;
DRAM[3424] = 8'b01010001;
DRAM[3425] = 8'b01111000;
DRAM[3426] = 8'b10001001;
DRAM[3427] = 8'b10010010;
DRAM[3428] = 8'b10001100;
DRAM[3429] = 8'b10001010;
DRAM[3430] = 8'b10010001;
DRAM[3431] = 8'b10010101;
DRAM[3432] = 8'b10010010;
DRAM[3433] = 8'b01000001;
DRAM[3434] = 8'b00101101;
DRAM[3435] = 8'b00101100;
DRAM[3436] = 8'b00101110;
DRAM[3437] = 8'b00110101;
DRAM[3438] = 8'b00110111;
DRAM[3439] = 8'b00110100;
DRAM[3440] = 8'b00110011;
DRAM[3441] = 8'b00101110;
DRAM[3442] = 8'b00111000;
DRAM[3443] = 8'b00101111;
DRAM[3444] = 8'b00110010;
DRAM[3445] = 8'b00110010;
DRAM[3446] = 8'b00110001;
DRAM[3447] = 8'b00111100;
DRAM[3448] = 8'b01101100;
DRAM[3449] = 8'b10010101;
DRAM[3450] = 8'b10001110;
DRAM[3451] = 8'b10001001;
DRAM[3452] = 8'b10011001;
DRAM[3453] = 8'b10100011;
DRAM[3454] = 8'b10100011;
DRAM[3455] = 8'b10100100;
DRAM[3456] = 8'b01011010;
DRAM[3457] = 8'b01011101;
DRAM[3458] = 8'b01011100;
DRAM[3459] = 8'b01011011;
DRAM[3460] = 8'b01011001;
DRAM[3461] = 8'b01010111;
DRAM[3462] = 8'b01101100;
DRAM[3463] = 8'b10001001;
DRAM[3464] = 8'b10011010;
DRAM[3465] = 8'b10100010;
DRAM[3466] = 8'b10100101;
DRAM[3467] = 8'b10100010;
DRAM[3468] = 8'b10100101;
DRAM[3469] = 8'b10011100;
DRAM[3470] = 8'b10000110;
DRAM[3471] = 8'b01101010;
DRAM[3472] = 8'b01001101;
DRAM[3473] = 8'b01010000;
DRAM[3474] = 8'b01010111;
DRAM[3475] = 8'b01011110;
DRAM[3476] = 8'b01100100;
DRAM[3477] = 8'b01100001;
DRAM[3478] = 8'b01100101;
DRAM[3479] = 8'b01100110;
DRAM[3480] = 8'b01100100;
DRAM[3481] = 8'b01100111;
DRAM[3482] = 8'b01101100;
DRAM[3483] = 8'b01101110;
DRAM[3484] = 8'b01110000;
DRAM[3485] = 8'b01110001;
DRAM[3486] = 8'b01110000;
DRAM[3487] = 8'b01101110;
DRAM[3488] = 8'b10101010;
DRAM[3489] = 8'b01110010;
DRAM[3490] = 8'b01100110;
DRAM[3491] = 8'b01101010;
DRAM[3492] = 8'b01110001;
DRAM[3493] = 8'b01101111;
DRAM[3494] = 8'b01110000;
DRAM[3495] = 8'b01110001;
DRAM[3496] = 8'b01111001;
DRAM[3497] = 8'b01111011;
DRAM[3498] = 8'b01111011;
DRAM[3499] = 8'b01111110;
DRAM[3500] = 8'b10000001;
DRAM[3501] = 8'b10001011;
DRAM[3502] = 8'b10000111;
DRAM[3503] = 8'b10000011;
DRAM[3504] = 8'b10001001;
DRAM[3505] = 8'b10001001;
DRAM[3506] = 8'b10001010;
DRAM[3507] = 8'b10000011;
DRAM[3508] = 8'b01111100;
DRAM[3509] = 8'b01110110;
DRAM[3510] = 8'b10000110;
DRAM[3511] = 8'b10101110;
DRAM[3512] = 8'b10111101;
DRAM[3513] = 8'b10111110;
DRAM[3514] = 8'b10111101;
DRAM[3515] = 8'b10111011;
DRAM[3516] = 8'b11000000;
DRAM[3517] = 8'b10111010;
DRAM[3518] = 8'b10111101;
DRAM[3519] = 8'b10111111;
DRAM[3520] = 8'b11000011;
DRAM[3521] = 8'b11000111;
DRAM[3522] = 8'b11001010;
DRAM[3523] = 8'b11001100;
DRAM[3524] = 8'b11001010;
DRAM[3525] = 8'b11001101;
DRAM[3526] = 8'b11001011;
DRAM[3527] = 8'b11001101;
DRAM[3528] = 8'b11001100;
DRAM[3529] = 8'b11001011;
DRAM[3530] = 8'b11001100;
DRAM[3531] = 8'b11001011;
DRAM[3532] = 8'b11001110;
DRAM[3533] = 8'b11010101;
DRAM[3534] = 8'b11011000;
DRAM[3535] = 8'b11100000;
DRAM[3536] = 8'b11000010;
DRAM[3537] = 8'b01001010;
DRAM[3538] = 8'b01010000;
DRAM[3539] = 8'b01110110;
DRAM[3540] = 8'b10001011;
DRAM[3541] = 8'b10010111;
DRAM[3542] = 8'b10011010;
DRAM[3543] = 8'b10011100;
DRAM[3544] = 8'b10011001;
DRAM[3545] = 8'b10010110;
DRAM[3546] = 8'b10000110;
DRAM[3547] = 8'b01100111;
DRAM[3548] = 8'b00111100;
DRAM[3549] = 8'b00101111;
DRAM[3550] = 8'b00101011;
DRAM[3551] = 8'b00101000;
DRAM[3552] = 8'b00110011;
DRAM[3553] = 8'b01011000;
DRAM[3554] = 8'b01110100;
DRAM[3555] = 8'b10100010;
DRAM[3556] = 8'b10101011;
DRAM[3557] = 8'b10010000;
DRAM[3558] = 8'b10010011;
DRAM[3559] = 8'b10010100;
DRAM[3560] = 8'b01100100;
DRAM[3561] = 8'b00101101;
DRAM[3562] = 8'b00101110;
DRAM[3563] = 8'b00101101;
DRAM[3564] = 8'b00110101;
DRAM[3565] = 8'b00110110;
DRAM[3566] = 8'b00110011;
DRAM[3567] = 8'b00110111;
DRAM[3568] = 8'b00110000;
DRAM[3569] = 8'b00110011;
DRAM[3570] = 8'b00110100;
DRAM[3571] = 8'b00110011;
DRAM[3572] = 8'b00111001;
DRAM[3573] = 8'b00101111;
DRAM[3574] = 8'b00101010;
DRAM[3575] = 8'b01011111;
DRAM[3576] = 8'b10010000;
DRAM[3577] = 8'b10010100;
DRAM[3578] = 8'b10001001;
DRAM[3579] = 8'b10010111;
DRAM[3580] = 8'b10011111;
DRAM[3581] = 8'b10100011;
DRAM[3582] = 8'b10100010;
DRAM[3583] = 8'b10100011;
DRAM[3584] = 8'b01011100;
DRAM[3585] = 8'b01011100;
DRAM[3586] = 8'b01011000;
DRAM[3587] = 8'b01011011;
DRAM[3588] = 8'b01010111;
DRAM[3589] = 8'b01010011;
DRAM[3590] = 8'b01101011;
DRAM[3591] = 8'b10001011;
DRAM[3592] = 8'b10011001;
DRAM[3593] = 8'b10100001;
DRAM[3594] = 8'b10100100;
DRAM[3595] = 8'b10100010;
DRAM[3596] = 8'b10100001;
DRAM[3597] = 8'b10011100;
DRAM[3598] = 8'b10001000;
DRAM[3599] = 8'b01101110;
DRAM[3600] = 8'b01001110;
DRAM[3601] = 8'b01010000;
DRAM[3602] = 8'b01011001;
DRAM[3603] = 8'b01011110;
DRAM[3604] = 8'b01011110;
DRAM[3605] = 8'b01100010;
DRAM[3606] = 8'b01100000;
DRAM[3607] = 8'b01100011;
DRAM[3608] = 8'b01100101;
DRAM[3609] = 8'b01101000;
DRAM[3610] = 8'b01101010;
DRAM[3611] = 8'b01101110;
DRAM[3612] = 8'b01110011;
DRAM[3613] = 8'b01110010;
DRAM[3614] = 8'b01101100;
DRAM[3615] = 8'b01110101;
DRAM[3616] = 8'b10111110;
DRAM[3617] = 8'b01101001;
DRAM[3618] = 8'b01101011;
DRAM[3619] = 8'b01100111;
DRAM[3620] = 8'b01101101;
DRAM[3621] = 8'b01110000;
DRAM[3622] = 8'b01110000;
DRAM[3623] = 8'b01101110;
DRAM[3624] = 8'b01110101;
DRAM[3625] = 8'b01110110;
DRAM[3626] = 8'b01111111;
DRAM[3627] = 8'b10000101;
DRAM[3628] = 8'b10000110;
DRAM[3629] = 8'b10000111;
DRAM[3630] = 8'b10001011;
DRAM[3631] = 8'b10000101;
DRAM[3632] = 8'b10001010;
DRAM[3633] = 8'b10001011;
DRAM[3634] = 8'b01111010;
DRAM[3635] = 8'b01111011;
DRAM[3636] = 8'b01110001;
DRAM[3637] = 8'b10010010;
DRAM[3638] = 8'b10110100;
DRAM[3639] = 8'b10111110;
DRAM[3640] = 8'b10111000;
DRAM[3641] = 8'b10111011;
DRAM[3642] = 8'b10111101;
DRAM[3643] = 8'b10111000;
DRAM[3644] = 8'b10101110;
DRAM[3645] = 8'b10111010;
DRAM[3646] = 8'b11000011;
DRAM[3647] = 8'b11000111;
DRAM[3648] = 8'b11000101;
DRAM[3649] = 8'b11000010;
DRAM[3650] = 8'b11001001;
DRAM[3651] = 8'b11001010;
DRAM[3652] = 8'b11001011;
DRAM[3653] = 8'b11001010;
DRAM[3654] = 8'b11001001;
DRAM[3655] = 8'b11001000;
DRAM[3656] = 8'b11001010;
DRAM[3657] = 8'b11001011;
DRAM[3658] = 8'b11010000;
DRAM[3659] = 8'b11010010;
DRAM[3660] = 8'b11001101;
DRAM[3661] = 8'b11010010;
DRAM[3662] = 8'b11010100;
DRAM[3663] = 8'b11011101;
DRAM[3664] = 8'b11100001;
DRAM[3665] = 8'b10000010;
DRAM[3666] = 8'b01001010;
DRAM[3667] = 8'b01110011;
DRAM[3668] = 8'b10001100;
DRAM[3669] = 8'b10010111;
DRAM[3670] = 8'b10010111;
DRAM[3671] = 8'b10011010;
DRAM[3672] = 8'b10011010;
DRAM[3673] = 8'b10011001;
DRAM[3674] = 8'b10000101;
DRAM[3675] = 8'b01101001;
DRAM[3676] = 8'b00111100;
DRAM[3677] = 8'b00101100;
DRAM[3678] = 8'b00101110;
DRAM[3679] = 8'b00100110;
DRAM[3680] = 8'b00100110;
DRAM[3681] = 8'b01011000;
DRAM[3682] = 8'b11001000;
DRAM[3683] = 8'b11010110;
DRAM[3684] = 8'b11001010;
DRAM[3685] = 8'b11001010;
DRAM[3686] = 8'b11010011;
DRAM[3687] = 8'b10101010;
DRAM[3688] = 8'b00101110;
DRAM[3689] = 8'b00101011;
DRAM[3690] = 8'b00101110;
DRAM[3691] = 8'b00101110;
DRAM[3692] = 8'b00110111;
DRAM[3693] = 8'b00110110;
DRAM[3694] = 8'b00111000;
DRAM[3695] = 8'b00110110;
DRAM[3696] = 8'b00110111;
DRAM[3697] = 8'b00110010;
DRAM[3698] = 8'b00101110;
DRAM[3699] = 8'b00110110;
DRAM[3700] = 8'b00101111;
DRAM[3701] = 8'b00101101;
DRAM[3702] = 8'b01001110;
DRAM[3703] = 8'b10001001;
DRAM[3704] = 8'b10010101;
DRAM[3705] = 8'b10001001;
DRAM[3706] = 8'b10010100;
DRAM[3707] = 8'b10100001;
DRAM[3708] = 8'b10100001;
DRAM[3709] = 8'b10011110;
DRAM[3710] = 8'b10011110;
DRAM[3711] = 8'b10011110;
DRAM[3712] = 8'b01011001;
DRAM[3713] = 8'b01011000;
DRAM[3714] = 8'b01011000;
DRAM[3715] = 8'b01011100;
DRAM[3716] = 8'b01011010;
DRAM[3717] = 8'b01010011;
DRAM[3718] = 8'b01101010;
DRAM[3719] = 8'b10000111;
DRAM[3720] = 8'b10011010;
DRAM[3721] = 8'b10100100;
DRAM[3722] = 8'b10100011;
DRAM[3723] = 8'b10100011;
DRAM[3724] = 8'b10100100;
DRAM[3725] = 8'b10011011;
DRAM[3726] = 8'b10001000;
DRAM[3727] = 8'b01101001;
DRAM[3728] = 8'b01001011;
DRAM[3729] = 8'b01001101;
DRAM[3730] = 8'b01010110;
DRAM[3731] = 8'b01010110;
DRAM[3732] = 8'b01011110;
DRAM[3733] = 8'b01100000;
DRAM[3734] = 8'b01011111;
DRAM[3735] = 8'b01011110;
DRAM[3736] = 8'b01100000;
DRAM[3737] = 8'b01101000;
DRAM[3738] = 8'b01101001;
DRAM[3739] = 8'b01101011;
DRAM[3740] = 8'b01101101;
DRAM[3741] = 8'b01101111;
DRAM[3742] = 8'b01100110;
DRAM[3743] = 8'b10100011;
DRAM[3744] = 8'b10101000;
DRAM[3745] = 8'b01101000;
DRAM[3746] = 8'b01100110;
DRAM[3747] = 8'b01101100;
DRAM[3748] = 8'b01101110;
DRAM[3749] = 8'b01110010;
DRAM[3750] = 8'b01110011;
DRAM[3751] = 8'b01110101;
DRAM[3752] = 8'b01110111;
DRAM[3753] = 8'b01111000;
DRAM[3754] = 8'b01111110;
DRAM[3755] = 8'b10000101;
DRAM[3756] = 8'b10001001;
DRAM[3757] = 8'b10000001;
DRAM[3758] = 8'b10000100;
DRAM[3759] = 8'b10000101;
DRAM[3760] = 8'b10001001;
DRAM[3761] = 8'b01111010;
DRAM[3762] = 8'b01110000;
DRAM[3763] = 8'b01111101;
DRAM[3764] = 8'b10011110;
DRAM[3765] = 8'b10110010;
DRAM[3766] = 8'b10110110;
DRAM[3767] = 8'b10110111;
DRAM[3768] = 8'b10110010;
DRAM[3769] = 8'b10110000;
DRAM[3770] = 8'b10110001;
DRAM[3771] = 8'b10111001;
DRAM[3772] = 8'b10111100;
DRAM[3773] = 8'b10111000;
DRAM[3774] = 8'b11000010;
DRAM[3775] = 8'b11000011;
DRAM[3776] = 8'b11000011;
DRAM[3777] = 8'b11000011;
DRAM[3778] = 8'b11000001;
DRAM[3779] = 8'b11000100;
DRAM[3780] = 8'b11000101;
DRAM[3781] = 8'b11000011;
DRAM[3782] = 8'b11000111;
DRAM[3783] = 8'b11001101;
DRAM[3784] = 8'b11001011;
DRAM[3785] = 8'b11001011;
DRAM[3786] = 8'b11001011;
DRAM[3787] = 8'b11001110;
DRAM[3788] = 8'b11010000;
DRAM[3789] = 8'b11001111;
DRAM[3790] = 8'b11010001;
DRAM[3791] = 8'b11010101;
DRAM[3792] = 8'b11100000;
DRAM[3793] = 8'b10111111;
DRAM[3794] = 8'b01000010;
DRAM[3795] = 8'b01101010;
DRAM[3796] = 8'b10001100;
DRAM[3797] = 8'b10010110;
DRAM[3798] = 8'b10011001;
DRAM[3799] = 8'b10011001;
DRAM[3800] = 8'b10011001;
DRAM[3801] = 8'b10010111;
DRAM[3802] = 8'b10000110;
DRAM[3803] = 8'b01100110;
DRAM[3804] = 8'b00111100;
DRAM[3805] = 8'b00101100;
DRAM[3806] = 8'b00100110;
DRAM[3807] = 8'b00100011;
DRAM[3808] = 8'b01101001;
DRAM[3809] = 8'b11011000;
DRAM[3810] = 8'b11001001;
DRAM[3811] = 8'b11000101;
DRAM[3812] = 8'b11010111;
DRAM[3813] = 8'b11100000;
DRAM[3814] = 8'b11100100;
DRAM[3815] = 8'b11011110;
DRAM[3816] = 8'b00101000;
DRAM[3817] = 8'b00101000;
DRAM[3818] = 8'b00101111;
DRAM[3819] = 8'b00111000;
DRAM[3820] = 8'b00110110;
DRAM[3821] = 8'b00110111;
DRAM[3822] = 8'b00110100;
DRAM[3823] = 8'b00110011;
DRAM[3824] = 8'b00110100;
DRAM[3825] = 8'b00110011;
DRAM[3826] = 8'b00110110;
DRAM[3827] = 8'b00111001;
DRAM[3828] = 8'b00101110;
DRAM[3829] = 8'b00110011;
DRAM[3830] = 8'b01111100;
DRAM[3831] = 8'b10010110;
DRAM[3832] = 8'b10001110;
DRAM[3833] = 8'b10001111;
DRAM[3834] = 8'b10011111;
DRAM[3835] = 8'b10100100;
DRAM[3836] = 8'b10100000;
DRAM[3837] = 8'b10011111;
DRAM[3838] = 8'b10011110;
DRAM[3839] = 8'b10011101;
DRAM[3840] = 8'b01011000;
DRAM[3841] = 8'b01011100;
DRAM[3842] = 8'b01011100;
DRAM[3843] = 8'b01011111;
DRAM[3844] = 8'b01011011;
DRAM[3845] = 8'b01011000;
DRAM[3846] = 8'b01101011;
DRAM[3847] = 8'b10001000;
DRAM[3848] = 8'b10011000;
DRAM[3849] = 8'b10100011;
DRAM[3850] = 8'b10100111;
DRAM[3851] = 8'b10100011;
DRAM[3852] = 8'b10100011;
DRAM[3853] = 8'b10011011;
DRAM[3854] = 8'b10001000;
DRAM[3855] = 8'b01100110;
DRAM[3856] = 8'b01001010;
DRAM[3857] = 8'b01001010;
DRAM[3858] = 8'b01010010;
DRAM[3859] = 8'b01011101;
DRAM[3860] = 8'b01100000;
DRAM[3861] = 8'b01100000;
DRAM[3862] = 8'b01100011;
DRAM[3863] = 8'b01100011;
DRAM[3864] = 8'b01100010;
DRAM[3865] = 8'b01100100;
DRAM[3866] = 8'b01101000;
DRAM[3867] = 8'b01101001;
DRAM[3868] = 8'b01101110;
DRAM[3869] = 8'b01110001;
DRAM[3870] = 8'b01100111;
DRAM[3871] = 8'b11001000;
DRAM[3872] = 8'b10100110;
DRAM[3873] = 8'b01101010;
DRAM[3874] = 8'b01100100;
DRAM[3875] = 8'b01101101;
DRAM[3876] = 8'b01101010;
DRAM[3877] = 8'b01110110;
DRAM[3878] = 8'b01110001;
DRAM[3879] = 8'b01110111;
DRAM[3880] = 8'b01110101;
DRAM[3881] = 8'b10000000;
DRAM[3882] = 8'b10000010;
DRAM[3883] = 8'b01111011;
DRAM[3884] = 8'b01110111;
DRAM[3885] = 8'b01111001;
DRAM[3886] = 8'b10000111;
DRAM[3887] = 8'b10000010;
DRAM[3888] = 8'b01111010;
DRAM[3889] = 8'b01101111;
DRAM[3890] = 8'b10000100;
DRAM[3891] = 8'b10100010;
DRAM[3892] = 8'b10110010;
DRAM[3893] = 8'b10110100;
DRAM[3894] = 8'b10100010;
DRAM[3895] = 8'b10101100;
DRAM[3896] = 8'b10110100;
DRAM[3897] = 8'b10101101;
DRAM[3898] = 8'b10110010;
DRAM[3899] = 8'b10110010;
DRAM[3900] = 8'b10111100;
DRAM[3901] = 8'b10111100;
DRAM[3902] = 8'b10111111;
DRAM[3903] = 8'b10111111;
DRAM[3904] = 8'b11000010;
DRAM[3905] = 8'b11000010;
DRAM[3906] = 8'b10111110;
DRAM[3907] = 8'b10111011;
DRAM[3908] = 8'b11000101;
DRAM[3909] = 8'b11001001;
DRAM[3910] = 8'b11001001;
DRAM[3911] = 8'b11001100;
DRAM[3912] = 8'b11001000;
DRAM[3913] = 8'b11000111;
DRAM[3914] = 8'b11000111;
DRAM[3915] = 8'b11001001;
DRAM[3916] = 8'b11001110;
DRAM[3917] = 8'b11001100;
DRAM[3918] = 8'b11001101;
DRAM[3919] = 8'b11001111;
DRAM[3920] = 8'b11011001;
DRAM[3921] = 8'b11011110;
DRAM[3922] = 8'b01110111;
DRAM[3923] = 8'b01100010;
DRAM[3924] = 8'b10000111;
DRAM[3925] = 8'b10011001;
DRAM[3926] = 8'b10011010;
DRAM[3927] = 8'b10011100;
DRAM[3928] = 8'b10011010;
DRAM[3929] = 8'b10010101;
DRAM[3930] = 8'b10000101;
DRAM[3931] = 8'b01100100;
DRAM[3932] = 8'b00110101;
DRAM[3933] = 8'b00100111;
DRAM[3934] = 8'b00101010;
DRAM[3935] = 8'b10011010;
DRAM[3936] = 8'b11010100;
DRAM[3937] = 8'b10110011;
DRAM[3938] = 8'b11001011;
DRAM[3939] = 8'b11011010;
DRAM[3940] = 8'b11011011;
DRAM[3941] = 8'b11011010;
DRAM[3942] = 8'b11011110;
DRAM[3943] = 8'b11101000;
DRAM[3944] = 8'b01110101;
DRAM[3945] = 8'b00101001;
DRAM[3946] = 8'b00101111;
DRAM[3947] = 8'b00110110;
DRAM[3948] = 8'b00110110;
DRAM[3949] = 8'b00110101;
DRAM[3950] = 8'b00110000;
DRAM[3951] = 8'b00110011;
DRAM[3952] = 8'b00101110;
DRAM[3953] = 8'b00101111;
DRAM[3954] = 8'b00111000;
DRAM[3955] = 8'b00110110;
DRAM[3956] = 8'b00110011;
DRAM[3957] = 8'b01101011;
DRAM[3958] = 8'b10010101;
DRAM[3959] = 8'b10010011;
DRAM[3960] = 8'b10001110;
DRAM[3961] = 8'b10011100;
DRAM[3962] = 8'b10011111;
DRAM[3963] = 8'b10100001;
DRAM[3964] = 8'b10011111;
DRAM[3965] = 8'b10011101;
DRAM[3966] = 8'b10011110;
DRAM[3967] = 8'b10011101;
DRAM[3968] = 8'b01011101;
DRAM[3969] = 8'b01011101;
DRAM[3970] = 8'b01011100;
DRAM[3971] = 8'b01100000;
DRAM[3972] = 8'b01011110;
DRAM[3973] = 8'b01011010;
DRAM[3974] = 8'b01101001;
DRAM[3975] = 8'b10000111;
DRAM[3976] = 8'b10010111;
DRAM[3977] = 8'b10100111;
DRAM[3978] = 8'b10100101;
DRAM[3979] = 8'b10100111;
DRAM[3980] = 8'b10100101;
DRAM[3981] = 8'b10011010;
DRAM[3982] = 8'b10001000;
DRAM[3983] = 8'b01100111;
DRAM[3984] = 8'b01001010;
DRAM[3985] = 8'b01001100;
DRAM[3986] = 8'b01010010;
DRAM[3987] = 8'b01011110;
DRAM[3988] = 8'b01100100;
DRAM[3989] = 8'b01100110;
DRAM[3990] = 8'b01100101;
DRAM[3991] = 8'b01100011;
DRAM[3992] = 8'b01100100;
DRAM[3993] = 8'b01100110;
DRAM[3994] = 8'b01101001;
DRAM[3995] = 8'b01101101;
DRAM[3996] = 8'b01110000;
DRAM[3997] = 8'b01110001;
DRAM[3998] = 8'b01101000;
DRAM[3999] = 8'b11010001;
DRAM[4000] = 8'b10010010;
DRAM[4001] = 8'b01011111;
DRAM[4002] = 8'b01100110;
DRAM[4003] = 8'b01100111;
DRAM[4004] = 8'b01101110;
DRAM[4005] = 8'b01101011;
DRAM[4006] = 8'b01101110;
DRAM[4007] = 8'b01110101;
DRAM[4008] = 8'b10000000;
DRAM[4009] = 8'b10000000;
DRAM[4010] = 8'b01111001;
DRAM[4011] = 8'b01110111;
DRAM[4012] = 8'b10000001;
DRAM[4013] = 8'b10000100;
DRAM[4014] = 8'b01111110;
DRAM[4015] = 8'b01111100;
DRAM[4016] = 8'b01101101;
DRAM[4017] = 8'b10000110;
DRAM[4018] = 8'b10101010;
DRAM[4019] = 8'b10110011;
DRAM[4020] = 8'b10101001;
DRAM[4021] = 8'b10100010;
DRAM[4022] = 8'b10101011;
DRAM[4023] = 8'b10101010;
DRAM[4024] = 8'b10110010;
DRAM[4025] = 8'b10110101;
DRAM[4026] = 8'b10110011;
DRAM[4027] = 8'b10110100;
DRAM[4028] = 8'b10111110;
DRAM[4029] = 8'b10111110;
DRAM[4030] = 8'b10111000;
DRAM[4031] = 8'b10111001;
DRAM[4032] = 8'b10111011;
DRAM[4033] = 8'b10111000;
DRAM[4034] = 8'b11000001;
DRAM[4035] = 8'b11000111;
DRAM[4036] = 8'b11000011;
DRAM[4037] = 8'b11000110;
DRAM[4038] = 8'b10111111;
DRAM[4039] = 8'b11001010;
DRAM[4040] = 8'b11000110;
DRAM[4041] = 8'b11001010;
DRAM[4042] = 8'b11001011;
DRAM[4043] = 8'b11001100;
DRAM[4044] = 8'b11001110;
DRAM[4045] = 8'b11001100;
DRAM[4046] = 8'b11001100;
DRAM[4047] = 8'b11001110;
DRAM[4048] = 8'b11010001;
DRAM[4049] = 8'b11010110;
DRAM[4050] = 8'b11010001;
DRAM[4051] = 8'b01100010;
DRAM[4052] = 8'b10000100;
DRAM[4053] = 8'b10010111;
DRAM[4054] = 8'b10011010;
DRAM[4055] = 8'b10011011;
DRAM[4056] = 8'b10011100;
DRAM[4057] = 8'b10010011;
DRAM[4058] = 8'b10000000;
DRAM[4059] = 8'b01011000;
DRAM[4060] = 8'b00101000;
DRAM[4061] = 8'b00111100;
DRAM[4062] = 8'b10110100;
DRAM[4063] = 8'b11000111;
DRAM[4064] = 8'b10101111;
DRAM[4065] = 8'b11010010;
DRAM[4066] = 8'b11011001;
DRAM[4067] = 8'b11010011;
DRAM[4068] = 8'b11010011;
DRAM[4069] = 8'b11001110;
DRAM[4070] = 8'b11010010;
DRAM[4071] = 8'b11100011;
DRAM[4072] = 8'b01111001;
DRAM[4073] = 8'b00101000;
DRAM[4074] = 8'b00101110;
DRAM[4075] = 8'b00110001;
DRAM[4076] = 8'b00110010;
DRAM[4077] = 8'b00101110;
DRAM[4078] = 8'b00110001;
DRAM[4079] = 8'b00101101;
DRAM[4080] = 8'b00101011;
DRAM[4081] = 8'b00110010;
DRAM[4082] = 8'b00111000;
DRAM[4083] = 8'b00101110;
DRAM[4084] = 8'b01001001;
DRAM[4085] = 8'b10010001;
DRAM[4086] = 8'b10011000;
DRAM[4087] = 8'b10001110;
DRAM[4088] = 8'b10011000;
DRAM[4089] = 8'b10011111;
DRAM[4090] = 8'b10011110;
DRAM[4091] = 8'b10011011;
DRAM[4092] = 8'b10011111;
DRAM[4093] = 8'b10011100;
DRAM[4094] = 8'b10011101;
DRAM[4095] = 8'b10011111;
DRAM[4096] = 8'b01011111;
DRAM[4097] = 8'b01100000;
DRAM[4098] = 8'b01100000;
DRAM[4099] = 8'b01100010;
DRAM[4100] = 8'b01100010;
DRAM[4101] = 8'b01011101;
DRAM[4102] = 8'b01101100;
DRAM[4103] = 8'b10001000;
DRAM[4104] = 8'b10011001;
DRAM[4105] = 8'b10100110;
DRAM[4106] = 8'b10100110;
DRAM[4107] = 8'b10100111;
DRAM[4108] = 8'b10100110;
DRAM[4109] = 8'b10011110;
DRAM[4110] = 8'b10001011;
DRAM[4111] = 8'b01101010;
DRAM[4112] = 8'b01001111;
DRAM[4113] = 8'b01010000;
DRAM[4114] = 8'b01011000;
DRAM[4115] = 8'b01011100;
DRAM[4116] = 8'b01100010;
DRAM[4117] = 8'b01100100;
DRAM[4118] = 8'b01100100;
DRAM[4119] = 8'b01100100;
DRAM[4120] = 8'b01100101;
DRAM[4121] = 8'b01101010;
DRAM[4122] = 8'b01101010;
DRAM[4123] = 8'b01101110;
DRAM[4124] = 8'b01110000;
DRAM[4125] = 8'b01101111;
DRAM[4126] = 8'b10000101;
DRAM[4127] = 8'b11001100;
DRAM[4128] = 8'b10010100;
DRAM[4129] = 8'b01100100;
DRAM[4130] = 8'b01100110;
DRAM[4131] = 8'b01101000;
DRAM[4132] = 8'b01100100;
DRAM[4133] = 8'b01110001;
DRAM[4134] = 8'b01110010;
DRAM[4135] = 8'b01111101;
DRAM[4136] = 8'b01111100;
DRAM[4137] = 8'b01110110;
DRAM[4138] = 8'b01111001;
DRAM[4139] = 8'b01111011;
DRAM[4140] = 8'b10000010;
DRAM[4141] = 8'b10000111;
DRAM[4142] = 8'b10000100;
DRAM[4143] = 8'b01101100;
DRAM[4144] = 8'b10000111;
DRAM[4145] = 8'b10100110;
DRAM[4146] = 8'b10100101;
DRAM[4147] = 8'b10100010;
DRAM[4148] = 8'b10101000;
DRAM[4149] = 8'b10100100;
DRAM[4150] = 8'b10100110;
DRAM[4151] = 8'b10110111;
DRAM[4152] = 8'b10110011;
DRAM[4153] = 8'b10101111;
DRAM[4154] = 8'b10111000;
DRAM[4155] = 8'b10111011;
DRAM[4156] = 8'b10110111;
DRAM[4157] = 8'b10111000;
DRAM[4158] = 8'b10111010;
DRAM[4159] = 8'b10101101;
DRAM[4160] = 8'b10110010;
DRAM[4161] = 8'b10111110;
DRAM[4162] = 8'b11000000;
DRAM[4163] = 8'b11000110;
DRAM[4164] = 8'b11000011;
DRAM[4165] = 8'b11000011;
DRAM[4166] = 8'b11000101;
DRAM[4167] = 8'b11000100;
DRAM[4168] = 8'b11001010;
DRAM[4169] = 8'b11000101;
DRAM[4170] = 8'b11000001;
DRAM[4171] = 8'b11000000;
DRAM[4172] = 8'b11000011;
DRAM[4173] = 8'b11001011;
DRAM[4174] = 8'b11001100;
DRAM[4175] = 8'b11001011;
DRAM[4176] = 8'b11001101;
DRAM[4177] = 8'b11001110;
DRAM[4178] = 8'b11010111;
DRAM[4179] = 8'b10111010;
DRAM[4180] = 8'b10000110;
DRAM[4181] = 8'b10010110;
DRAM[4182] = 8'b10011000;
DRAM[4183] = 8'b10011101;
DRAM[4184] = 8'b10011010;
DRAM[4185] = 8'b10010001;
DRAM[4186] = 8'b01110101;
DRAM[4187] = 8'b01001110;
DRAM[4188] = 8'b01111000;
DRAM[4189] = 8'b11001111;
DRAM[4190] = 8'b11000001;
DRAM[4191] = 8'b10111001;
DRAM[4192] = 8'b11010100;
DRAM[4193] = 8'b11010100;
DRAM[4194] = 8'b11010001;
DRAM[4195] = 8'b11001011;
DRAM[4196] = 8'b11001011;
DRAM[4197] = 8'b11001111;
DRAM[4198] = 8'b11011001;
DRAM[4199] = 8'b11100100;
DRAM[4200] = 8'b01111001;
DRAM[4201] = 8'b00100111;
DRAM[4202] = 8'b00110101;
DRAM[4203] = 8'b00110110;
DRAM[4204] = 8'b00110000;
DRAM[4205] = 8'b00101100;
DRAM[4206] = 8'b00101110;
DRAM[4207] = 8'b00101100;
DRAM[4208] = 8'b00110011;
DRAM[4209] = 8'b00110011;
DRAM[4210] = 8'b00100110;
DRAM[4211] = 8'b00110011;
DRAM[4212] = 8'b01111011;
DRAM[4213] = 8'b10011001;
DRAM[4214] = 8'b10010010;
DRAM[4215] = 8'b10010111;
DRAM[4216] = 8'b10100001;
DRAM[4217] = 8'b10011110;
DRAM[4218] = 8'b10011110;
DRAM[4219] = 8'b10011101;
DRAM[4220] = 8'b10011110;
DRAM[4221] = 8'b10011100;
DRAM[4222] = 8'b10011010;
DRAM[4223] = 8'b10011101;
DRAM[4224] = 8'b01100010;
DRAM[4225] = 8'b01100101;
DRAM[4226] = 8'b01100011;
DRAM[4227] = 8'b01100101;
DRAM[4228] = 8'b01100000;
DRAM[4229] = 8'b01011110;
DRAM[4230] = 8'b01101011;
DRAM[4231] = 8'b10000111;
DRAM[4232] = 8'b10011001;
DRAM[4233] = 8'b10100100;
DRAM[4234] = 8'b10101000;
DRAM[4235] = 8'b10100111;
DRAM[4236] = 8'b10101010;
DRAM[4237] = 8'b10100000;
DRAM[4238] = 8'b10001000;
DRAM[4239] = 8'b01101010;
DRAM[4240] = 8'b01010000;
DRAM[4241] = 8'b01001111;
DRAM[4242] = 8'b01011000;
DRAM[4243] = 8'b01011111;
DRAM[4244] = 8'b01100100;
DRAM[4245] = 8'b01100110;
DRAM[4246] = 8'b01100111;
DRAM[4247] = 8'b01100110;
DRAM[4248] = 8'b01100101;
DRAM[4249] = 8'b01101000;
DRAM[4250] = 8'b01101111;
DRAM[4251] = 8'b01101110;
DRAM[4252] = 8'b01110010;
DRAM[4253] = 8'b01101100;
DRAM[4254] = 8'b10100001;
DRAM[4255] = 8'b11001001;
DRAM[4256] = 8'b01111101;
DRAM[4257] = 8'b01100111;
DRAM[4258] = 8'b01011110;
DRAM[4259] = 8'b01100111;
DRAM[4260] = 8'b01101111;
DRAM[4261] = 8'b01101111;
DRAM[4262] = 8'b01101101;
DRAM[4263] = 8'b01110111;
DRAM[4264] = 8'b01110011;
DRAM[4265] = 8'b01111010;
DRAM[4266] = 8'b01111101;
DRAM[4267] = 8'b10000001;
DRAM[4268] = 8'b01110111;
DRAM[4269] = 8'b01111000;
DRAM[4270] = 8'b01101000;
DRAM[4271] = 8'b10001010;
DRAM[4272] = 8'b10100001;
DRAM[4273] = 8'b10011010;
DRAM[4274] = 8'b10011000;
DRAM[4275] = 8'b10011010;
DRAM[4276] = 8'b10100001;
DRAM[4277] = 8'b10100111;
DRAM[4278] = 8'b10101011;
DRAM[4279] = 8'b10110000;
DRAM[4280] = 8'b10110100;
DRAM[4281] = 8'b10111000;
DRAM[4282] = 8'b10101100;
DRAM[4283] = 8'b10110101;
DRAM[4284] = 8'b10110011;
DRAM[4285] = 8'b10110011;
DRAM[4286] = 8'b10101000;
DRAM[4287] = 8'b10110011;
DRAM[4288] = 8'b10110111;
DRAM[4289] = 8'b10111100;
DRAM[4290] = 8'b10110111;
DRAM[4291] = 8'b10111110;
DRAM[4292] = 8'b11000010;
DRAM[4293] = 8'b11000011;
DRAM[4294] = 8'b11000111;
DRAM[4295] = 8'b11000101;
DRAM[4296] = 8'b11000111;
DRAM[4297] = 8'b10110101;
DRAM[4298] = 8'b10101110;
DRAM[4299] = 8'b11000100;
DRAM[4300] = 8'b11001000;
DRAM[4301] = 8'b11001010;
DRAM[4302] = 8'b11001001;
DRAM[4303] = 8'b11001001;
DRAM[4304] = 8'b11000111;
DRAM[4305] = 8'b11001001;
DRAM[4306] = 8'b11001110;
DRAM[4307] = 8'b11010100;
DRAM[4308] = 8'b11000100;
DRAM[4309] = 8'b10010010;
DRAM[4310] = 8'b10011001;
DRAM[4311] = 8'b10010111;
DRAM[4312] = 8'b10010100;
DRAM[4313] = 8'b10001001;
DRAM[4314] = 8'b01111111;
DRAM[4315] = 8'b10110110;
DRAM[4316] = 8'b11001100;
DRAM[4317] = 8'b10111100;
DRAM[4318] = 8'b11000101;
DRAM[4319] = 8'b11010100;
DRAM[4320] = 8'b11010010;
DRAM[4321] = 8'b11001100;
DRAM[4322] = 8'b11001010;
DRAM[4323] = 8'b11001001;
DRAM[4324] = 8'b11001101;
DRAM[4325] = 8'b11010011;
DRAM[4326] = 8'b11011010;
DRAM[4327] = 8'b11011111;
DRAM[4328] = 8'b01111010;
DRAM[4329] = 8'b00101011;
DRAM[4330] = 8'b00110000;
DRAM[4331] = 8'b00110011;
DRAM[4332] = 8'b00110011;
DRAM[4333] = 8'b00110010;
DRAM[4334] = 8'b00110000;
DRAM[4335] = 8'b00110101;
DRAM[4336] = 8'b00110110;
DRAM[4337] = 8'b00110010;
DRAM[4338] = 8'b00100001;
DRAM[4339] = 8'b01011001;
DRAM[4340] = 8'b10010101;
DRAM[4341] = 8'b10010110;
DRAM[4342] = 8'b10010001;
DRAM[4343] = 8'b10011111;
DRAM[4344] = 8'b10011110;
DRAM[4345] = 8'b10011101;
DRAM[4346] = 8'b10011100;
DRAM[4347] = 8'b10011100;
DRAM[4348] = 8'b10011011;
DRAM[4349] = 8'b10011100;
DRAM[4350] = 8'b10011010;
DRAM[4351] = 8'b10011010;
DRAM[4352] = 8'b01100011;
DRAM[4353] = 8'b01100110;
DRAM[4354] = 8'b01100110;
DRAM[4355] = 8'b01100011;
DRAM[4356] = 8'b01100011;
DRAM[4357] = 8'b01100100;
DRAM[4358] = 8'b01110001;
DRAM[4359] = 8'b10001000;
DRAM[4360] = 8'b10011010;
DRAM[4361] = 8'b10100001;
DRAM[4362] = 8'b10100110;
DRAM[4363] = 8'b10101100;
DRAM[4364] = 8'b10101000;
DRAM[4365] = 8'b10100000;
DRAM[4366] = 8'b10001100;
DRAM[4367] = 8'b01101101;
DRAM[4368] = 8'b01001110;
DRAM[4369] = 8'b01010001;
DRAM[4370] = 8'b01011010;
DRAM[4371] = 8'b01100000;
DRAM[4372] = 8'b01100100;
DRAM[4373] = 8'b01100101;
DRAM[4374] = 8'b01100111;
DRAM[4375] = 8'b01100100;
DRAM[4376] = 8'b01100101;
DRAM[4377] = 8'b01100101;
DRAM[4378] = 8'b01101011;
DRAM[4379] = 8'b01101011;
DRAM[4380] = 8'b01101101;
DRAM[4381] = 8'b01100100;
DRAM[4382] = 8'b10100100;
DRAM[4383] = 8'b10110100;
DRAM[4384] = 8'b10000010;
DRAM[4385] = 8'b01101100;
DRAM[4386] = 8'b01100101;
DRAM[4387] = 8'b01101001;
DRAM[4388] = 8'b01100110;
DRAM[4389] = 8'b01100110;
DRAM[4390] = 8'b01101111;
DRAM[4391] = 8'b01110100;
DRAM[4392] = 8'b01110011;
DRAM[4393] = 8'b01111101;
DRAM[4394] = 8'b01111110;
DRAM[4395] = 8'b01110100;
DRAM[4396] = 8'b01111001;
DRAM[4397] = 8'b01110010;
DRAM[4398] = 8'b10001001;
DRAM[4399] = 8'b10011101;
DRAM[4400] = 8'b10011001;
DRAM[4401] = 8'b10010011;
DRAM[4402] = 8'b10010001;
DRAM[4403] = 8'b10010110;
DRAM[4404] = 8'b10011110;
DRAM[4405] = 8'b10101010;
DRAM[4406] = 8'b10110010;
DRAM[4407] = 8'b10110010;
DRAM[4408] = 8'b10100111;
DRAM[4409] = 8'b10101001;
DRAM[4410] = 8'b10110110;
DRAM[4411] = 8'b10110011;
DRAM[4412] = 8'b10101110;
DRAM[4413] = 8'b10100111;
DRAM[4414] = 8'b10110001;
DRAM[4415] = 8'b10110111;
DRAM[4416] = 8'b10111000;
DRAM[4417] = 8'b10110111;
DRAM[4418] = 8'b10111000;
DRAM[4419] = 8'b10110111;
DRAM[4420] = 8'b10111011;
DRAM[4421] = 8'b10111111;
DRAM[4422] = 8'b11000101;
DRAM[4423] = 8'b11001001;
DRAM[4424] = 8'b10110100;
DRAM[4425] = 8'b10110010;
DRAM[4426] = 8'b10111110;
DRAM[4427] = 8'b11000010;
DRAM[4428] = 8'b11000101;
DRAM[4429] = 8'b11000110;
DRAM[4430] = 8'b11000101;
DRAM[4431] = 8'b11000110;
DRAM[4432] = 8'b11000110;
DRAM[4433] = 8'b11000100;
DRAM[4434] = 8'b11000011;
DRAM[4435] = 8'b11000111;
DRAM[4436] = 8'b11010001;
DRAM[4437] = 8'b10101000;
DRAM[4438] = 8'b10010111;
DRAM[4439] = 8'b10010010;
DRAM[4440] = 8'b10010001;
DRAM[4441] = 8'b10111001;
DRAM[4442] = 8'b11001111;
DRAM[4443] = 8'b11000000;
DRAM[4444] = 8'b10111100;
DRAM[4445] = 8'b11001001;
DRAM[4446] = 8'b11010010;
DRAM[4447] = 8'b11001110;
DRAM[4448] = 8'b11001010;
DRAM[4449] = 8'b11001010;
DRAM[4450] = 8'b11001010;
DRAM[4451] = 8'b11001011;
DRAM[4452] = 8'b11010010;
DRAM[4453] = 8'b11010110;
DRAM[4454] = 8'b11011100;
DRAM[4455] = 8'b11011111;
DRAM[4456] = 8'b01010011;
DRAM[4457] = 8'b00101101;
DRAM[4458] = 8'b00110110;
DRAM[4459] = 8'b00110001;
DRAM[4460] = 8'b00110001;
DRAM[4461] = 8'b00101110;
DRAM[4462] = 8'b00101010;
DRAM[4463] = 8'b00110000;
DRAM[4464] = 8'b00110101;
DRAM[4465] = 8'b00101110;
DRAM[4466] = 8'b01000000;
DRAM[4467] = 8'b10000111;
DRAM[4468] = 8'b10011010;
DRAM[4469] = 8'b10010001;
DRAM[4470] = 8'b10011010;
DRAM[4471] = 8'b10100001;
DRAM[4472] = 8'b10011111;
DRAM[4473] = 8'b10011110;
DRAM[4474] = 8'b10011101;
DRAM[4475] = 8'b10011100;
DRAM[4476] = 8'b10011100;
DRAM[4477] = 8'b10011100;
DRAM[4478] = 8'b10011000;
DRAM[4479] = 8'b10011011;
DRAM[4480] = 8'b01100101;
DRAM[4481] = 8'b01100001;
DRAM[4482] = 8'b01100000;
DRAM[4483] = 8'b01100011;
DRAM[4484] = 8'b01100110;
DRAM[4485] = 8'b01100011;
DRAM[4486] = 8'b01110010;
DRAM[4487] = 8'b10001001;
DRAM[4488] = 8'b10011100;
DRAM[4489] = 8'b10100101;
DRAM[4490] = 8'b10101011;
DRAM[4491] = 8'b10101100;
DRAM[4492] = 8'b10101100;
DRAM[4493] = 8'b10100101;
DRAM[4494] = 8'b10001101;
DRAM[4495] = 8'b01101010;
DRAM[4496] = 8'b01001100;
DRAM[4497] = 8'b01010010;
DRAM[4498] = 8'b01011100;
DRAM[4499] = 8'b01100001;
DRAM[4500] = 8'b01100100;
DRAM[4501] = 8'b01100101;
DRAM[4502] = 8'b01100101;
DRAM[4503] = 8'b01100110;
DRAM[4504] = 8'b01100100;
DRAM[4505] = 8'b01100101;
DRAM[4506] = 8'b01101011;
DRAM[4507] = 8'b01101100;
DRAM[4508] = 8'b01100111;
DRAM[4509] = 8'b01011110;
DRAM[4510] = 8'b11001011;
DRAM[4511] = 8'b10101110;
DRAM[4512] = 8'b10000011;
DRAM[4513] = 8'b01101101;
DRAM[4514] = 8'b01101000;
DRAM[4515] = 8'b01101010;
DRAM[4516] = 8'b01101001;
DRAM[4517] = 8'b01101010;
DRAM[4518] = 8'b01101100;
DRAM[4519] = 8'b01101110;
DRAM[4520] = 8'b01111010;
DRAM[4521] = 8'b01110011;
DRAM[4522] = 8'b01110110;
DRAM[4523] = 8'b01111100;
DRAM[4524] = 8'b01110100;
DRAM[4525] = 8'b10010001;
DRAM[4526] = 8'b10010101;
DRAM[4527] = 8'b10010001;
DRAM[4528] = 8'b10001110;
DRAM[4529] = 8'b10010011;
DRAM[4530] = 8'b10000111;
DRAM[4531] = 8'b10100000;
DRAM[4532] = 8'b10100010;
DRAM[4533] = 8'b10100110;
DRAM[4534] = 8'b10101100;
DRAM[4535] = 8'b10101010;
DRAM[4536] = 8'b10100100;
DRAM[4537] = 8'b10110000;
DRAM[4538] = 8'b10110001;
DRAM[4539] = 8'b10101010;
DRAM[4540] = 8'b10100001;
DRAM[4541] = 8'b10110100;
DRAM[4542] = 8'b10101101;
DRAM[4543] = 8'b10101111;
DRAM[4544] = 8'b10110011;
DRAM[4545] = 8'b10110000;
DRAM[4546] = 8'b10110011;
DRAM[4547] = 8'b10110100;
DRAM[4548] = 8'b10110110;
DRAM[4549] = 8'b10111010;
DRAM[4550] = 8'b10101101;
DRAM[4551] = 8'b10110000;
DRAM[4552] = 8'b10111001;
DRAM[4553] = 8'b10110011;
DRAM[4554] = 8'b10110111;
DRAM[4555] = 8'b10111001;
DRAM[4556] = 8'b11000001;
DRAM[4557] = 8'b11000100;
DRAM[4558] = 8'b11000000;
DRAM[4559] = 8'b10111101;
DRAM[4560] = 8'b10111110;
DRAM[4561] = 8'b11000011;
DRAM[4562] = 8'b10111100;
DRAM[4563] = 8'b10111100;
DRAM[4564] = 8'b11000010;
DRAM[4565] = 8'b10111001;
DRAM[4566] = 8'b10010100;
DRAM[4567] = 8'b10100110;
DRAM[4568] = 8'b11001010;
DRAM[4569] = 8'b11001001;
DRAM[4570] = 8'b10111101;
DRAM[4571] = 8'b11000001;
DRAM[4572] = 8'b11010001;
DRAM[4573] = 8'b11001110;
DRAM[4574] = 8'b11001001;
DRAM[4575] = 8'b11001000;
DRAM[4576] = 8'b11001001;
DRAM[4577] = 8'b11001100;
DRAM[4578] = 8'b11001100;
DRAM[4579] = 8'b11001011;
DRAM[4580] = 8'b11010000;
DRAM[4581] = 8'b11010101;
DRAM[4582] = 8'b11011100;
DRAM[4583] = 8'b11100001;
DRAM[4584] = 8'b00101010;
DRAM[4585] = 8'b00101111;
DRAM[4586] = 8'b00110101;
DRAM[4587] = 8'b00110011;
DRAM[4588] = 8'b00110000;
DRAM[4589] = 8'b00101010;
DRAM[4590] = 8'b00110000;
DRAM[4591] = 8'b00110100;
DRAM[4592] = 8'b00111000;
DRAM[4593] = 8'b00111110;
DRAM[4594] = 8'b01101011;
DRAM[4595] = 8'b10010101;
DRAM[4596] = 8'b10010011;
DRAM[4597] = 8'b10010110;
DRAM[4598] = 8'b10100000;
DRAM[4599] = 8'b10011111;
DRAM[4600] = 8'b10011101;
DRAM[4601] = 8'b10011101;
DRAM[4602] = 8'b10011101;
DRAM[4603] = 8'b10011110;
DRAM[4604] = 8'b10011001;
DRAM[4605] = 8'b10011011;
DRAM[4606] = 8'b10011001;
DRAM[4607] = 8'b10011001;
DRAM[4608] = 8'b01100100;
DRAM[4609] = 8'b01100101;
DRAM[4610] = 8'b01100010;
DRAM[4611] = 8'b01100010;
DRAM[4612] = 8'b01100100;
DRAM[4613] = 8'b01100100;
DRAM[4614] = 8'b01110001;
DRAM[4615] = 8'b10001010;
DRAM[4616] = 8'b10011101;
DRAM[4617] = 8'b10101000;
DRAM[4618] = 8'b10101010;
DRAM[4619] = 8'b10101011;
DRAM[4620] = 8'b10101101;
DRAM[4621] = 8'b10100110;
DRAM[4622] = 8'b10001110;
DRAM[4623] = 8'b01101100;
DRAM[4624] = 8'b01001111;
DRAM[4625] = 8'b01001110;
DRAM[4626] = 8'b01011000;
DRAM[4627] = 8'b01011100;
DRAM[4628] = 8'b01100011;
DRAM[4629] = 8'b01100110;
DRAM[4630] = 8'b01100001;
DRAM[4631] = 8'b01100001;
DRAM[4632] = 8'b01100100;
DRAM[4633] = 8'b01100010;
DRAM[4634] = 8'b01100101;
DRAM[4635] = 8'b01101001;
DRAM[4636] = 8'b01100100;
DRAM[4637] = 8'b01011000;
DRAM[4638] = 8'b11011000;
DRAM[4639] = 8'b10110000;
DRAM[4640] = 8'b10001011;
DRAM[4641] = 8'b01110110;
DRAM[4642] = 8'b01100101;
DRAM[4643] = 8'b01101010;
DRAM[4644] = 8'b01100110;
DRAM[4645] = 8'b01101110;
DRAM[4646] = 8'b01110001;
DRAM[4647] = 8'b01110001;
DRAM[4648] = 8'b01110110;
DRAM[4649] = 8'b01110111;
DRAM[4650] = 8'b01111010;
DRAM[4651] = 8'b01110010;
DRAM[4652] = 8'b10001010;
DRAM[4653] = 8'b10010010;
DRAM[4654] = 8'b10010110;
DRAM[4655] = 8'b10001011;
DRAM[4656] = 8'b10001101;
DRAM[4657] = 8'b10000100;
DRAM[4658] = 8'b10010110;
DRAM[4659] = 8'b10011110;
DRAM[4660] = 8'b10100011;
DRAM[4661] = 8'b10011110;
DRAM[4662] = 8'b10011111;
DRAM[4663] = 8'b10101101;
DRAM[4664] = 8'b10110100;
DRAM[4665] = 8'b10100110;
DRAM[4666] = 8'b10011110;
DRAM[4667] = 8'b10101010;
DRAM[4668] = 8'b10110000;
DRAM[4669] = 8'b10101011;
DRAM[4670] = 8'b10110000;
DRAM[4671] = 8'b10101100;
DRAM[4672] = 8'b10101111;
DRAM[4673] = 8'b10101110;
DRAM[4674] = 8'b10110010;
DRAM[4675] = 8'b10111111;
DRAM[4676] = 8'b10111001;
DRAM[4677] = 8'b10110011;
DRAM[4678] = 8'b10110101;
DRAM[4679] = 8'b10111001;
DRAM[4680] = 8'b10111100;
DRAM[4681] = 8'b10110111;
DRAM[4682] = 8'b10111111;
DRAM[4683] = 8'b10111110;
DRAM[4684] = 8'b10111111;
DRAM[4685] = 8'b10111010;
DRAM[4686] = 8'b10111000;
DRAM[4687] = 8'b10111001;
DRAM[4688] = 8'b10111100;
DRAM[4689] = 8'b10111000;
DRAM[4690] = 8'b10110100;
DRAM[4691] = 8'b10110111;
DRAM[4692] = 8'b10111000;
DRAM[4693] = 8'b11000000;
DRAM[4694] = 8'b10111110;
DRAM[4695] = 8'b11001001;
DRAM[4696] = 8'b10111101;
DRAM[4697] = 8'b11000000;
DRAM[4698] = 8'b11001110;
DRAM[4699] = 8'b11001101;
DRAM[4700] = 8'b11001100;
DRAM[4701] = 8'b11001001;
DRAM[4702] = 8'b11000110;
DRAM[4703] = 8'b11001001;
DRAM[4704] = 8'b11001100;
DRAM[4705] = 8'b11001100;
DRAM[4706] = 8'b11001100;
DRAM[4707] = 8'b11000110;
DRAM[4708] = 8'b11010000;
DRAM[4709] = 8'b11010100;
DRAM[4710] = 8'b11011110;
DRAM[4711] = 8'b11011001;
DRAM[4712] = 8'b00100000;
DRAM[4713] = 8'b00101111;
DRAM[4714] = 8'b00110000;
DRAM[4715] = 8'b00110001;
DRAM[4716] = 8'b00110011;
DRAM[4717] = 8'b00101010;
DRAM[4718] = 8'b00110100;
DRAM[4719] = 8'b00110100;
DRAM[4720] = 8'b01000000;
DRAM[4721] = 8'b01011010;
DRAM[4722] = 8'b10010000;
DRAM[4723] = 8'b10010101;
DRAM[4724] = 8'b10010010;
DRAM[4725] = 8'b10011100;
DRAM[4726] = 8'b10100001;
DRAM[4727] = 8'b10100000;
DRAM[4728] = 8'b10100000;
DRAM[4729] = 8'b10011100;
DRAM[4730] = 8'b10011100;
DRAM[4731] = 8'b10011101;
DRAM[4732] = 8'b10011010;
DRAM[4733] = 8'b10011011;
DRAM[4734] = 8'b10011010;
DRAM[4735] = 8'b10011100;
DRAM[4736] = 8'b01100100;
DRAM[4737] = 8'b01100011;
DRAM[4738] = 8'b01100010;
DRAM[4739] = 8'b01100000;
DRAM[4740] = 8'b01100010;
DRAM[4741] = 8'b01100101;
DRAM[4742] = 8'b01110000;
DRAM[4743] = 8'b10001010;
DRAM[4744] = 8'b10011101;
DRAM[4745] = 8'b10101001;
DRAM[4746] = 8'b10101101;
DRAM[4747] = 8'b10101110;
DRAM[4748] = 8'b10101100;
DRAM[4749] = 8'b10100100;
DRAM[4750] = 8'b10001100;
DRAM[4751] = 8'b01101010;
DRAM[4752] = 8'b01001101;
DRAM[4753] = 8'b01001110;
DRAM[4754] = 8'b01010111;
DRAM[4755] = 8'b01011110;
DRAM[4756] = 8'b01100001;
DRAM[4757] = 8'b01100010;
DRAM[4758] = 8'b01100011;
DRAM[4759] = 8'b01100001;
DRAM[4760] = 8'b01100010;
DRAM[4761] = 8'b01100111;
DRAM[4762] = 8'b01100111;
DRAM[4763] = 8'b01101010;
DRAM[4764] = 8'b01100100;
DRAM[4765] = 8'b01100010;
DRAM[4766] = 8'b11010100;
DRAM[4767] = 8'b10110001;
DRAM[4768] = 8'b10010100;
DRAM[4769] = 8'b10000001;
DRAM[4770] = 8'b01111000;
DRAM[4771] = 8'b01101110;
DRAM[4772] = 8'b01101011;
DRAM[4773] = 8'b01101100;
DRAM[4774] = 8'b01101101;
DRAM[4775] = 8'b01101111;
DRAM[4776] = 8'b01110111;
DRAM[4777] = 8'b01111011;
DRAM[4778] = 8'b01110011;
DRAM[4779] = 8'b10000111;
DRAM[4780] = 8'b10010100;
DRAM[4781] = 8'b10001101;
DRAM[4782] = 8'b10001110;
DRAM[4783] = 8'b10010001;
DRAM[4784] = 8'b10001000;
DRAM[4785] = 8'b10010100;
DRAM[4786] = 8'b10010111;
DRAM[4787] = 8'b10010100;
DRAM[4788] = 8'b10011000;
DRAM[4789] = 8'b10011101;
DRAM[4790] = 8'b10101101;
DRAM[4791] = 8'b10101010;
DRAM[4792] = 8'b10100011;
DRAM[4793] = 8'b10011110;
DRAM[4794] = 8'b10101100;
DRAM[4795] = 8'b10101011;
DRAM[4796] = 8'b10101010;
DRAM[4797] = 8'b10110000;
DRAM[4798] = 8'b10101101;
DRAM[4799] = 8'b10101110;
DRAM[4800] = 8'b10101111;
DRAM[4801] = 8'b10101010;
DRAM[4802] = 8'b10101100;
DRAM[4803] = 8'b10110000;
DRAM[4804] = 8'b10110110;
DRAM[4805] = 8'b10111001;
DRAM[4806] = 8'b10110110;
DRAM[4807] = 8'b10110000;
DRAM[4808] = 8'b10110111;
DRAM[4809] = 8'b10111111;
DRAM[4810] = 8'b10111010;
DRAM[4811] = 8'b10111100;
DRAM[4812] = 8'b10110101;
DRAM[4813] = 8'b10110000;
DRAM[4814] = 8'b10101111;
DRAM[4815] = 8'b10111001;
DRAM[4816] = 8'b10110101;
DRAM[4817] = 8'b10110000;
DRAM[4818] = 8'b10101100;
DRAM[4819] = 8'b10100111;
DRAM[4820] = 8'b11000001;
DRAM[4821] = 8'b10111110;
DRAM[4822] = 8'b10111000;
DRAM[4823] = 8'b11000011;
DRAM[4824] = 8'b11000111;
DRAM[4825] = 8'b11010001;
DRAM[4826] = 8'b11001101;
DRAM[4827] = 8'b11000100;
DRAM[4828] = 8'b11001000;
DRAM[4829] = 8'b11001000;
DRAM[4830] = 8'b11000111;
DRAM[4831] = 8'b11001001;
DRAM[4832] = 8'b11001011;
DRAM[4833] = 8'b11001101;
DRAM[4834] = 8'b10111111;
DRAM[4835] = 8'b10111011;
DRAM[4836] = 8'b11001011;
DRAM[4837] = 8'b11010001;
DRAM[4838] = 8'b11011011;
DRAM[4839] = 8'b10010000;
DRAM[4840] = 8'b00100110;
DRAM[4841] = 8'b00101111;
DRAM[4842] = 8'b00101111;
DRAM[4843] = 8'b00110101;
DRAM[4844] = 8'b00101101;
DRAM[4845] = 8'b00101100;
DRAM[4846] = 8'b00110111;
DRAM[4847] = 8'b00110100;
DRAM[4848] = 8'b01000001;
DRAM[4849] = 8'b10000000;
DRAM[4850] = 8'b10010110;
DRAM[4851] = 8'b10010000;
DRAM[4852] = 8'b10010111;
DRAM[4853] = 8'b10011111;
DRAM[4854] = 8'b10100010;
DRAM[4855] = 8'b10100000;
DRAM[4856] = 8'b10011111;
DRAM[4857] = 8'b10011100;
DRAM[4858] = 8'b10011110;
DRAM[4859] = 8'b10011110;
DRAM[4860] = 8'b10011100;
DRAM[4861] = 8'b10011011;
DRAM[4862] = 8'b10011100;
DRAM[4863] = 8'b10011100;
DRAM[4864] = 8'b01100001;
DRAM[4865] = 8'b01100101;
DRAM[4866] = 8'b01100100;
DRAM[4867] = 8'b01100010;
DRAM[4868] = 8'b01100000;
DRAM[4869] = 8'b01100001;
DRAM[4870] = 8'b01101101;
DRAM[4871] = 8'b10000111;
DRAM[4872] = 8'b10011011;
DRAM[4873] = 8'b10100111;
DRAM[4874] = 8'b10101100;
DRAM[4875] = 8'b10101101;
DRAM[4876] = 8'b10101100;
DRAM[4877] = 8'b10100101;
DRAM[4878] = 8'b10001111;
DRAM[4879] = 8'b01101101;
DRAM[4880] = 8'b01010010;
DRAM[4881] = 8'b01001111;
DRAM[4882] = 8'b01011010;
DRAM[4883] = 8'b01011110;
DRAM[4884] = 8'b01100010;
DRAM[4885] = 8'b01100011;
DRAM[4886] = 8'b01100010;
DRAM[4887] = 8'b01100011;
DRAM[4888] = 8'b01100100;
DRAM[4889] = 8'b01100011;
DRAM[4890] = 8'b01100111;
DRAM[4891] = 8'b01101010;
DRAM[4892] = 8'b01100011;
DRAM[4893] = 8'b01110101;
DRAM[4894] = 8'b11001111;
DRAM[4895] = 8'b10110000;
DRAM[4896] = 8'b10011001;
DRAM[4897] = 8'b10001110;
DRAM[4898] = 8'b01111110;
DRAM[4899] = 8'b01110001;
DRAM[4900] = 8'b01101001;
DRAM[4901] = 8'b01101000;
DRAM[4902] = 8'b01110001;
DRAM[4903] = 8'b01110100;
DRAM[4904] = 8'b01101111;
DRAM[4905] = 8'b01101011;
DRAM[4906] = 8'b10001010;
DRAM[4907] = 8'b10001110;
DRAM[4908] = 8'b10010000;
DRAM[4909] = 8'b10001100;
DRAM[4910] = 8'b10001010;
DRAM[4911] = 8'b10000011;
DRAM[4912] = 8'b10010100;
DRAM[4913] = 8'b10010100;
DRAM[4914] = 8'b10011001;
DRAM[4915] = 8'b10001001;
DRAM[4916] = 8'b10010101;
DRAM[4917] = 8'b10011110;
DRAM[4918] = 8'b10100001;
DRAM[4919] = 8'b10100011;
DRAM[4920] = 8'b10011011;
DRAM[4921] = 8'b10101110;
DRAM[4922] = 8'b10101100;
DRAM[4923] = 8'b10100110;
DRAM[4924] = 8'b10101000;
DRAM[4925] = 8'b10110000;
DRAM[4926] = 8'b10110000;
DRAM[4927] = 8'b10101110;
DRAM[4928] = 8'b10100101;
DRAM[4929] = 8'b10101100;
DRAM[4930] = 8'b10100101;
DRAM[4931] = 8'b10101100;
DRAM[4932] = 8'b10101111;
DRAM[4933] = 8'b10101001;
DRAM[4934] = 8'b10110100;
DRAM[4935] = 8'b10111010;
DRAM[4936] = 8'b10110011;
DRAM[4937] = 8'b10111011;
DRAM[4938] = 8'b10111001;
DRAM[4939] = 8'b10110010;
DRAM[4940] = 8'b10110110;
DRAM[4941] = 8'b10110111;
DRAM[4942] = 8'b10101111;
DRAM[4943] = 8'b10101100;
DRAM[4944] = 8'b10110001;
DRAM[4945] = 8'b10100010;
DRAM[4946] = 8'b10110001;
DRAM[4947] = 8'b11000010;
DRAM[4948] = 8'b10111010;
DRAM[4949] = 8'b10111001;
DRAM[4950] = 8'b11001000;
DRAM[4951] = 8'b11001101;
DRAM[4952] = 8'b11001011;
DRAM[4953] = 8'b11001010;
DRAM[4954] = 8'b11000101;
DRAM[4955] = 8'b11001000;
DRAM[4956] = 8'b11001000;
DRAM[4957] = 8'b11001000;
DRAM[4958] = 8'b11001000;
DRAM[4959] = 8'b11001100;
DRAM[4960] = 8'b11001100;
DRAM[4961] = 8'b11000100;
DRAM[4962] = 8'b10100010;
DRAM[4963] = 8'b10101010;
DRAM[4964] = 8'b11000001;
DRAM[4965] = 8'b11000111;
DRAM[4966] = 8'b11010101;
DRAM[4967] = 8'b01011100;
DRAM[4968] = 8'b00101010;
DRAM[4969] = 8'b00101111;
DRAM[4970] = 8'b00101111;
DRAM[4971] = 8'b00110100;
DRAM[4972] = 8'b00101100;
DRAM[4973] = 8'b00110001;
DRAM[4974] = 8'b00110011;
DRAM[4975] = 8'b00110010;
DRAM[4976] = 8'b01010100;
DRAM[4977] = 8'b10010100;
DRAM[4978] = 8'b10010101;
DRAM[4979] = 8'b10010101;
DRAM[4980] = 8'b10011111;
DRAM[4981] = 8'b10100001;
DRAM[4982] = 8'b10100000;
DRAM[4983] = 8'b10011111;
DRAM[4984] = 8'b10100001;
DRAM[4985] = 8'b10011110;
DRAM[4986] = 8'b10011100;
DRAM[4987] = 8'b10011110;
DRAM[4988] = 8'b10011101;
DRAM[4989] = 8'b10011101;
DRAM[4990] = 8'b10011100;
DRAM[4991] = 8'b10011100;
DRAM[4992] = 8'b01100010;
DRAM[4993] = 8'b01100011;
DRAM[4994] = 8'b01011110;
DRAM[4995] = 8'b01100000;
DRAM[4996] = 8'b01100001;
DRAM[4997] = 8'b01100010;
DRAM[4998] = 8'b01101110;
DRAM[4999] = 8'b10001100;
DRAM[5000] = 8'b10011111;
DRAM[5001] = 8'b10101010;
DRAM[5002] = 8'b10101011;
DRAM[5003] = 8'b10101101;
DRAM[5004] = 8'b10101000;
DRAM[5005] = 8'b10100010;
DRAM[5006] = 8'b10001101;
DRAM[5007] = 8'b01101010;
DRAM[5008] = 8'b01010010;
DRAM[5009] = 8'b01010000;
DRAM[5010] = 8'b01011010;
DRAM[5011] = 8'b01011110;
DRAM[5012] = 8'b01100100;
DRAM[5013] = 8'b01100100;
DRAM[5014] = 8'b01100011;
DRAM[5015] = 8'b01100011;
DRAM[5016] = 8'b01100010;
DRAM[5017] = 8'b01100101;
DRAM[5018] = 8'b01100101;
DRAM[5019] = 8'b01100101;
DRAM[5020] = 8'b01100011;
DRAM[5021] = 8'b01110110;
DRAM[5022] = 8'b11001010;
DRAM[5023] = 8'b10101110;
DRAM[5024] = 8'b10011111;
DRAM[5025] = 8'b10010000;
DRAM[5026] = 8'b10000101;
DRAM[5027] = 8'b10000000;
DRAM[5028] = 8'b01101000;
DRAM[5029] = 8'b01100010;
DRAM[5030] = 8'b01101011;
DRAM[5031] = 8'b01110100;
DRAM[5032] = 8'b01101110;
DRAM[5033] = 8'b10000101;
DRAM[5034] = 8'b10001100;
DRAM[5035] = 8'b10001001;
DRAM[5036] = 8'b10001110;
DRAM[5037] = 8'b10000000;
DRAM[5038] = 8'b01111011;
DRAM[5039] = 8'b10010011;
DRAM[5040] = 8'b10011000;
DRAM[5041] = 8'b10010001;
DRAM[5042] = 8'b10010000;
DRAM[5043] = 8'b10011000;
DRAM[5044] = 8'b10010110;
DRAM[5045] = 8'b10010000;
DRAM[5046] = 8'b10011000;
DRAM[5047] = 8'b10011100;
DRAM[5048] = 8'b10101011;
DRAM[5049] = 8'b10101001;
DRAM[5050] = 8'b10100011;
DRAM[5051] = 8'b10101001;
DRAM[5052] = 8'b10101010;
DRAM[5053] = 8'b10100011;
DRAM[5054] = 8'b10101010;
DRAM[5055] = 8'b10100001;
DRAM[5056] = 8'b10100110;
DRAM[5057] = 8'b10100100;
DRAM[5058] = 8'b10100101;
DRAM[5059] = 8'b10100000;
DRAM[5060] = 8'b10100111;
DRAM[5061] = 8'b10110000;
DRAM[5062] = 8'b10101100;
DRAM[5063] = 8'b10110000;
DRAM[5064] = 8'b10111000;
DRAM[5065] = 8'b10101110;
DRAM[5066] = 8'b10110001;
DRAM[5067] = 8'b10101101;
DRAM[5068] = 8'b10101010;
DRAM[5069] = 8'b10110101;
DRAM[5070] = 8'b10101001;
DRAM[5071] = 8'b10011100;
DRAM[5072] = 8'b10101010;
DRAM[5073] = 8'b10111111;
DRAM[5074] = 8'b10111011;
DRAM[5075] = 8'b10111011;
DRAM[5076] = 8'b11000100;
DRAM[5077] = 8'b11001010;
DRAM[5078] = 8'b11001000;
DRAM[5079] = 8'b11000110;
DRAM[5080] = 8'b11000000;
DRAM[5081] = 8'b11000000;
DRAM[5082] = 8'b11000101;
DRAM[5083] = 8'b11000111;
DRAM[5084] = 8'b11001010;
DRAM[5085] = 8'b11001000;
DRAM[5086] = 8'b11001011;
DRAM[5087] = 8'b11001101;
DRAM[5088] = 8'b11001101;
DRAM[5089] = 8'b10100110;
DRAM[5090] = 8'b10100000;
DRAM[5091] = 8'b10101010;
DRAM[5092] = 8'b10001110;
DRAM[5093] = 8'b10111011;
DRAM[5094] = 8'b11001011;
DRAM[5095] = 8'b00100100;
DRAM[5096] = 8'b00110000;
DRAM[5097] = 8'b00111001;
DRAM[5098] = 8'b00110110;
DRAM[5099] = 8'b00101100;
DRAM[5100] = 8'b00101100;
DRAM[5101] = 8'b00110000;
DRAM[5102] = 8'b00110010;
DRAM[5103] = 8'b01010100;
DRAM[5104] = 8'b10000001;
DRAM[5105] = 8'b10010101;
DRAM[5106] = 8'b10010000;
DRAM[5107] = 8'b10011011;
DRAM[5108] = 8'b10011110;
DRAM[5109] = 8'b10100000;
DRAM[5110] = 8'b10011110;
DRAM[5111] = 8'b10100000;
DRAM[5112] = 8'b10011110;
DRAM[5113] = 8'b10011101;
DRAM[5114] = 8'b10011101;
DRAM[5115] = 8'b10011100;
DRAM[5116] = 8'b10011110;
DRAM[5117] = 8'b10011110;
DRAM[5118] = 8'b10011100;
DRAM[5119] = 8'b10011110;
DRAM[5120] = 8'b01100011;
DRAM[5121] = 8'b01011101;
DRAM[5122] = 8'b01100000;
DRAM[5123] = 8'b01011101;
DRAM[5124] = 8'b01011110;
DRAM[5125] = 8'b01011111;
DRAM[5126] = 8'b01101111;
DRAM[5127] = 8'b10001011;
DRAM[5128] = 8'b10011101;
DRAM[5129] = 8'b10101000;
DRAM[5130] = 8'b10101100;
DRAM[5131] = 8'b10101011;
DRAM[5132] = 8'b10101010;
DRAM[5133] = 8'b10100011;
DRAM[5134] = 8'b10010000;
DRAM[5135] = 8'b01101111;
DRAM[5136] = 8'b01010010;
DRAM[5137] = 8'b01010010;
DRAM[5138] = 8'b01011011;
DRAM[5139] = 8'b01100000;
DRAM[5140] = 8'b01100010;
DRAM[5141] = 8'b01100011;
DRAM[5142] = 8'b01100011;
DRAM[5143] = 8'b01100000;
DRAM[5144] = 8'b01100010;
DRAM[5145] = 8'b01100011;
DRAM[5146] = 8'b01100100;
DRAM[5147] = 8'b01100010;
DRAM[5148] = 8'b01011100;
DRAM[5149] = 8'b10001100;
DRAM[5150] = 8'b11000001;
DRAM[5151] = 8'b10101100;
DRAM[5152] = 8'b10011110;
DRAM[5153] = 8'b10010010;
DRAM[5154] = 8'b10000111;
DRAM[5155] = 8'b10000010;
DRAM[5156] = 8'b01101000;
DRAM[5157] = 8'b01100100;
DRAM[5158] = 8'b01101011;
DRAM[5159] = 8'b01101010;
DRAM[5160] = 8'b10000111;
DRAM[5161] = 8'b10001001;
DRAM[5162] = 8'b10000100;
DRAM[5163] = 8'b10001011;
DRAM[5164] = 8'b01111101;
DRAM[5165] = 8'b01111100;
DRAM[5166] = 8'b10010000;
DRAM[5167] = 8'b10001101;
DRAM[5168] = 8'b10001110;
DRAM[5169] = 8'b10010000;
DRAM[5170] = 8'b10010000;
DRAM[5171] = 8'b10001010;
DRAM[5172] = 8'b10011011;
DRAM[5173] = 8'b10010100;
DRAM[5174] = 8'b10011001;
DRAM[5175] = 8'b10100011;
DRAM[5176] = 8'b10011011;
DRAM[5177] = 8'b10011111;
DRAM[5178] = 8'b10101011;
DRAM[5179] = 8'b10100001;
DRAM[5180] = 8'b10100001;
DRAM[5181] = 8'b10100011;
DRAM[5182] = 8'b10100001;
DRAM[5183] = 8'b10101001;
DRAM[5184] = 8'b10011111;
DRAM[5185] = 8'b10100000;
DRAM[5186] = 8'b10100010;
DRAM[5187] = 8'b10100110;
DRAM[5188] = 8'b10100111;
DRAM[5189] = 8'b10101100;
DRAM[5190] = 8'b10101100;
DRAM[5191] = 8'b10101001;
DRAM[5192] = 8'b10101100;
DRAM[5193] = 8'b10101100;
DRAM[5194] = 8'b10101000;
DRAM[5195] = 8'b10101100;
DRAM[5196] = 8'b10100110;
DRAM[5197] = 8'b10100010;
DRAM[5198] = 8'b10100100;
DRAM[5199] = 8'b10110100;
DRAM[5200] = 8'b10111010;
DRAM[5201] = 8'b10110011;
DRAM[5202] = 8'b10111111;
DRAM[5203] = 8'b11001011;
DRAM[5204] = 8'b11001011;
DRAM[5205] = 8'b11000101;
DRAM[5206] = 8'b11000000;
DRAM[5207] = 8'b11000000;
DRAM[5208] = 8'b11000010;
DRAM[5209] = 8'b11000101;
DRAM[5210] = 8'b11000110;
DRAM[5211] = 8'b11001010;
DRAM[5212] = 8'b11001000;
DRAM[5213] = 8'b11001010;
DRAM[5214] = 8'b11001110;
DRAM[5215] = 8'b11010000;
DRAM[5216] = 8'b10111100;
DRAM[5217] = 8'b10011110;
DRAM[5218] = 8'b10101000;
DRAM[5219] = 8'b10001101;
DRAM[5220] = 8'b10100011;
DRAM[5221] = 8'b10111100;
DRAM[5222] = 8'b01111111;
DRAM[5223] = 8'b00101000;
DRAM[5224] = 8'b00101011;
DRAM[5225] = 8'b00110111;
DRAM[5226] = 8'b00101101;
DRAM[5227] = 8'b00101001;
DRAM[5228] = 8'b00110011;
DRAM[5229] = 8'b00101111;
DRAM[5230] = 8'b00111111;
DRAM[5231] = 8'b01101001;
DRAM[5232] = 8'b10011000;
DRAM[5233] = 8'b10010010;
DRAM[5234] = 8'b10010011;
DRAM[5235] = 8'b10011110;
DRAM[5236] = 8'b10100000;
DRAM[5237] = 8'b10100001;
DRAM[5238] = 8'b10011110;
DRAM[5239] = 8'b10011110;
DRAM[5240] = 8'b10011111;
DRAM[5241] = 8'b10100000;
DRAM[5242] = 8'b10011110;
DRAM[5243] = 8'b10011100;
DRAM[5244] = 8'b10011100;
DRAM[5245] = 8'b10011110;
DRAM[5246] = 8'b10011110;
DRAM[5247] = 8'b10011111;
DRAM[5248] = 8'b01100000;
DRAM[5249] = 8'b01100000;
DRAM[5250] = 8'b01011100;
DRAM[5251] = 8'b01100000;
DRAM[5252] = 8'b01011100;
DRAM[5253] = 8'b01100001;
DRAM[5254] = 8'b01110010;
DRAM[5255] = 8'b10001101;
DRAM[5256] = 8'b10011110;
DRAM[5257] = 8'b10100111;
DRAM[5258] = 8'b10101100;
DRAM[5259] = 8'b10101010;
DRAM[5260] = 8'b10101100;
DRAM[5261] = 8'b10100101;
DRAM[5262] = 8'b10001110;
DRAM[5263] = 8'b01101110;
DRAM[5264] = 8'b01001110;
DRAM[5265] = 8'b01010100;
DRAM[5266] = 8'b01011011;
DRAM[5267] = 8'b01100001;
DRAM[5268] = 8'b01100100;
DRAM[5269] = 8'b01100001;
DRAM[5270] = 8'b01100011;
DRAM[5271] = 8'b01100010;
DRAM[5272] = 8'b01100001;
DRAM[5273] = 8'b01100010;
DRAM[5274] = 8'b01100011;
DRAM[5275] = 8'b01100001;
DRAM[5276] = 8'b01011001;
DRAM[5277] = 8'b10011010;
DRAM[5278] = 8'b11000000;
DRAM[5279] = 8'b10110110;
DRAM[5280] = 8'b10100001;
DRAM[5281] = 8'b10011101;
DRAM[5282] = 8'b10010000;
DRAM[5283] = 8'b10000111;
DRAM[5284] = 8'b01110011;
DRAM[5285] = 8'b01101011;
DRAM[5286] = 8'b01100100;
DRAM[5287] = 8'b10000011;
DRAM[5288] = 8'b10001100;
DRAM[5289] = 8'b10000111;
DRAM[5290] = 8'b10001010;
DRAM[5291] = 8'b01111000;
DRAM[5292] = 8'b01111100;
DRAM[5293] = 8'b10010010;
DRAM[5294] = 8'b10010001;
DRAM[5295] = 8'b10001110;
DRAM[5296] = 8'b10001011;
DRAM[5297] = 8'b01111111;
DRAM[5298] = 8'b10001110;
DRAM[5299] = 8'b10011000;
DRAM[5300] = 8'b10001100;
DRAM[5301] = 8'b10011000;
DRAM[5302] = 8'b10100001;
DRAM[5303] = 8'b10011001;
DRAM[5304] = 8'b10100000;
DRAM[5305] = 8'b10011010;
DRAM[5306] = 8'b10011011;
DRAM[5307] = 8'b10010100;
DRAM[5308] = 8'b10011101;
DRAM[5309] = 8'b10100101;
DRAM[5310] = 8'b10011111;
DRAM[5311] = 8'b10011001;
DRAM[5312] = 8'b10011101;
DRAM[5313] = 8'b10100110;
DRAM[5314] = 8'b10100011;
DRAM[5315] = 8'b10101000;
DRAM[5316] = 8'b10100011;
DRAM[5317] = 8'b10100110;
DRAM[5318] = 8'b10100101;
DRAM[5319] = 8'b10100110;
DRAM[5320] = 8'b10100001;
DRAM[5321] = 8'b10100000;
DRAM[5322] = 8'b10100110;
DRAM[5323] = 8'b10100001;
DRAM[5324] = 8'b10011000;
DRAM[5325] = 8'b10101011;
DRAM[5326] = 8'b10111001;
DRAM[5327] = 8'b10110000;
DRAM[5328] = 8'b10111011;
DRAM[5329] = 8'b11000101;
DRAM[5330] = 8'b11000101;
DRAM[5331] = 8'b11000000;
DRAM[5332] = 8'b10111101;
DRAM[5333] = 8'b10111110;
DRAM[5334] = 8'b11000010;
DRAM[5335] = 8'b11000101;
DRAM[5336] = 8'b11000101;
DRAM[5337] = 8'b11001000;
DRAM[5338] = 8'b11001011;
DRAM[5339] = 8'b11001001;
DRAM[5340] = 8'b11001010;
DRAM[5341] = 8'b11001110;
DRAM[5342] = 8'b11010001;
DRAM[5343] = 8'b11001111;
DRAM[5344] = 8'b10011000;
DRAM[5345] = 8'b10100100;
DRAM[5346] = 8'b10011001;
DRAM[5347] = 8'b10100001;
DRAM[5348] = 8'b10011010;
DRAM[5349] = 8'b11010101;
DRAM[5350] = 8'b01000010;
DRAM[5351] = 8'b00101100;
DRAM[5352] = 8'b00101111;
DRAM[5353] = 8'b00110001;
DRAM[5354] = 8'b00110010;
DRAM[5355] = 8'b00110101;
DRAM[5356] = 8'b00110011;
DRAM[5357] = 8'b00110111;
DRAM[5358] = 8'b01001110;
DRAM[5359] = 8'b10001110;
DRAM[5360] = 8'b10011001;
DRAM[5361] = 8'b10010000;
DRAM[5362] = 8'b10011010;
DRAM[5363] = 8'b10011110;
DRAM[5364] = 8'b10100000;
DRAM[5365] = 8'b10011101;
DRAM[5366] = 8'b10011110;
DRAM[5367] = 8'b10011110;
DRAM[5368] = 8'b10011110;
DRAM[5369] = 8'b10011101;
DRAM[5370] = 8'b10011100;
DRAM[5371] = 8'b10011100;
DRAM[5372] = 8'b10011110;
DRAM[5373] = 8'b10011011;
DRAM[5374] = 8'b10011100;
DRAM[5375] = 8'b10011101;
DRAM[5376] = 8'b01100000;
DRAM[5377] = 8'b01100000;
DRAM[5378] = 8'b01100000;
DRAM[5379] = 8'b01011110;
DRAM[5380] = 8'b01100010;
DRAM[5381] = 8'b01100101;
DRAM[5382] = 8'b01110100;
DRAM[5383] = 8'b10001100;
DRAM[5384] = 8'b10011110;
DRAM[5385] = 8'b10101000;
DRAM[5386] = 8'b10101011;
DRAM[5387] = 8'b10101110;
DRAM[5388] = 8'b10101011;
DRAM[5389] = 8'b10100100;
DRAM[5390] = 8'b10010010;
DRAM[5391] = 8'b01101100;
DRAM[5392] = 8'b01001110;
DRAM[5393] = 8'b01010000;
DRAM[5394] = 8'b01011001;
DRAM[5395] = 8'b01100000;
DRAM[5396] = 8'b01100001;
DRAM[5397] = 8'b01100000;
DRAM[5398] = 8'b01011100;
DRAM[5399] = 8'b01100010;
DRAM[5400] = 8'b01100010;
DRAM[5401] = 8'b01100010;
DRAM[5402] = 8'b01100100;
DRAM[5403] = 8'b01100000;
DRAM[5404] = 8'b01010110;
DRAM[5405] = 8'b10011010;
DRAM[5406] = 8'b11001010;
DRAM[5407] = 8'b11000001;
DRAM[5408] = 8'b10101111;
DRAM[5409] = 8'b10100111;
DRAM[5410] = 8'b10001101;
DRAM[5411] = 8'b10010010;
DRAM[5412] = 8'b01111101;
DRAM[5413] = 8'b01100000;
DRAM[5414] = 8'b01111100;
DRAM[5415] = 8'b10001000;
DRAM[5416] = 8'b10000000;
DRAM[5417] = 8'b10001001;
DRAM[5418] = 8'b01111000;
DRAM[5419] = 8'b01111111;
DRAM[5420] = 8'b10001111;
DRAM[5421] = 8'b10001001;
DRAM[5422] = 8'b10001101;
DRAM[5423] = 8'b10000111;
DRAM[5424] = 8'b01111111;
DRAM[5425] = 8'b10000111;
DRAM[5426] = 8'b10010111;
DRAM[5427] = 8'b10001001;
DRAM[5428] = 8'b10010000;
DRAM[5429] = 8'b10011110;
DRAM[5430] = 8'b10011001;
DRAM[5431] = 8'b10000000;
DRAM[5432] = 8'b01111111;
DRAM[5433] = 8'b10001101;
DRAM[5434] = 8'b10010111;
DRAM[5435] = 8'b10000111;
DRAM[5436] = 8'b10001000;
DRAM[5437] = 8'b01101010;
DRAM[5438] = 8'b01111011;
DRAM[5439] = 8'b10100010;
DRAM[5440] = 8'b10100100;
DRAM[5441] = 8'b10011110;
DRAM[5442] = 8'b10100000;
DRAM[5443] = 8'b10100001;
DRAM[5444] = 8'b10100101;
DRAM[5445] = 8'b10011110;
DRAM[5446] = 8'b10100001;
DRAM[5447] = 8'b10100010;
DRAM[5448] = 8'b10100010;
DRAM[5449] = 8'b10100000;
DRAM[5450] = 8'b10010100;
DRAM[5451] = 8'b10011110;
DRAM[5452] = 8'b10111100;
DRAM[5453] = 8'b10110000;
DRAM[5454] = 8'b10110001;
DRAM[5455] = 8'b11000001;
DRAM[5456] = 8'b11001001;
DRAM[5457] = 8'b11000010;
DRAM[5458] = 8'b10111100;
DRAM[5459] = 8'b10111100;
DRAM[5460] = 8'b10111111;
DRAM[5461] = 8'b11000011;
DRAM[5462] = 8'b11000010;
DRAM[5463] = 8'b11000101;
DRAM[5464] = 8'b11001001;
DRAM[5465] = 8'b11001011;
DRAM[5466] = 8'b11001011;
DRAM[5467] = 8'b11001100;
DRAM[5468] = 8'b11001101;
DRAM[5469] = 8'b11010001;
DRAM[5470] = 8'b11010010;
DRAM[5471] = 8'b10110010;
DRAM[5472] = 8'b10100001;
DRAM[5473] = 8'b10001111;
DRAM[5474] = 8'b01111100;
DRAM[5475] = 8'b01101100;
DRAM[5476] = 8'b10110110;
DRAM[5477] = 8'b11000010;
DRAM[5478] = 8'b00100100;
DRAM[5479] = 8'b00101100;
DRAM[5480] = 8'b00110000;
DRAM[5481] = 8'b00110100;
DRAM[5482] = 8'b00110011;
DRAM[5483] = 8'b00111100;
DRAM[5484] = 8'b00110111;
DRAM[5485] = 8'b00110111;
DRAM[5486] = 8'b01100111;
DRAM[5487] = 8'b10011000;
DRAM[5488] = 8'b10010001;
DRAM[5489] = 8'b10010110;
DRAM[5490] = 8'b10011110;
DRAM[5491] = 8'b10011111;
DRAM[5492] = 8'b10011101;
DRAM[5493] = 8'b10011101;
DRAM[5494] = 8'b10011011;
DRAM[5495] = 8'b10011011;
DRAM[5496] = 8'b10011111;
DRAM[5497] = 8'b10011100;
DRAM[5498] = 8'b10011011;
DRAM[5499] = 8'b10011100;
DRAM[5500] = 8'b10011101;
DRAM[5501] = 8'b10011101;
DRAM[5502] = 8'b10011101;
DRAM[5503] = 8'b10011011;
DRAM[5504] = 8'b01100010;
DRAM[5505] = 8'b01100011;
DRAM[5506] = 8'b01100000;
DRAM[5507] = 8'b01100011;
DRAM[5508] = 8'b01100100;
DRAM[5509] = 8'b01101001;
DRAM[5510] = 8'b01110101;
DRAM[5511] = 8'b10001110;
DRAM[5512] = 8'b10011101;
DRAM[5513] = 8'b10101100;
DRAM[5514] = 8'b10101100;
DRAM[5515] = 8'b10101101;
DRAM[5516] = 8'b10101101;
DRAM[5517] = 8'b10100110;
DRAM[5518] = 8'b10010101;
DRAM[5519] = 8'b01101100;
DRAM[5520] = 8'b01001010;
DRAM[5521] = 8'b01001100;
DRAM[5522] = 8'b01011000;
DRAM[5523] = 8'b01011110;
DRAM[5524] = 8'b01100001;
DRAM[5525] = 8'b01100010;
DRAM[5526] = 8'b01100100;
DRAM[5527] = 8'b01100010;
DRAM[5528] = 8'b01100100;
DRAM[5529] = 8'b01100100;
DRAM[5530] = 8'b01100010;
DRAM[5531] = 8'b01011111;
DRAM[5532] = 8'b01010100;
DRAM[5533] = 8'b10011001;
DRAM[5534] = 8'b11001101;
DRAM[5535] = 8'b11000011;
DRAM[5536] = 8'b10101110;
DRAM[5537] = 8'b10100001;
DRAM[5538] = 8'b10010110;
DRAM[5539] = 8'b10011000;
DRAM[5540] = 8'b10000110;
DRAM[5541] = 8'b01110101;
DRAM[5542] = 8'b01111010;
DRAM[5543] = 8'b10000000;
DRAM[5544] = 8'b10000101;
DRAM[5545] = 8'b01101110;
DRAM[5546] = 8'b01111100;
DRAM[5547] = 8'b10001011;
DRAM[5548] = 8'b10001100;
DRAM[5549] = 8'b10001000;
DRAM[5550] = 8'b10001000;
DRAM[5551] = 8'b01111100;
DRAM[5552] = 8'b10000111;
DRAM[5553] = 8'b10010001;
DRAM[5554] = 8'b10000101;
DRAM[5555] = 8'b10010001;
DRAM[5556] = 8'b10010111;
DRAM[5557] = 8'b10000000;
DRAM[5558] = 8'b01101111;
DRAM[5559] = 8'b10000111;
DRAM[5560] = 8'b01111000;
DRAM[5561] = 8'b01101010;
DRAM[5562] = 8'b01101001;
DRAM[5563] = 8'b01110011;
DRAM[5564] = 8'b10100000;
DRAM[5565] = 8'b10011110;
DRAM[5566] = 8'b01110110;
DRAM[5567] = 8'b01111110;
DRAM[5568] = 8'b10000001;
DRAM[5569] = 8'b10011100;
DRAM[5570] = 8'b10010110;
DRAM[5571] = 8'b10001111;
DRAM[5572] = 8'b10001010;
DRAM[5573] = 8'b10011001;
DRAM[5574] = 8'b10000111;
DRAM[5575] = 8'b01001110;
DRAM[5576] = 8'b10000001;
DRAM[5577] = 8'b10010011;
DRAM[5578] = 8'b10100000;
DRAM[5579] = 8'b10111000;
DRAM[5580] = 8'b10100111;
DRAM[5581] = 8'b10111001;
DRAM[5582] = 8'b11001001;
DRAM[5583] = 8'b11000101;
DRAM[5584] = 8'b11000011;
DRAM[5585] = 8'b11000000;
DRAM[5586] = 8'b11000000;
DRAM[5587] = 8'b11000000;
DRAM[5588] = 8'b11000010;
DRAM[5589] = 8'b11000110;
DRAM[5590] = 8'b11001000;
DRAM[5591] = 8'b11001001;
DRAM[5592] = 8'b11001100;
DRAM[5593] = 8'b11001101;
DRAM[5594] = 8'b11001100;
DRAM[5595] = 8'b11001100;
DRAM[5596] = 8'b11001110;
DRAM[5597] = 8'b11010010;
DRAM[5598] = 8'b11001000;
DRAM[5599] = 8'b10100011;
DRAM[5600] = 8'b01110010;
DRAM[5601] = 8'b01010110;
DRAM[5602] = 8'b01100010;
DRAM[5603] = 8'b10010101;
DRAM[5604] = 8'b11010110;
DRAM[5605] = 8'b01101011;
DRAM[5606] = 8'b00100101;
DRAM[5607] = 8'b00101000;
DRAM[5608] = 8'b00110011;
DRAM[5609] = 8'b00101101;
DRAM[5610] = 8'b00110001;
DRAM[5611] = 8'b00111000;
DRAM[5612] = 8'b00110100;
DRAM[5613] = 8'b01001000;
DRAM[5614] = 8'b10001100;
DRAM[5615] = 8'b10010110;
DRAM[5616] = 8'b10010010;
DRAM[5617] = 8'b10011100;
DRAM[5618] = 8'b10100000;
DRAM[5619] = 8'b10011101;
DRAM[5620] = 8'b10100000;
DRAM[5621] = 8'b10011101;
DRAM[5622] = 8'b10011100;
DRAM[5623] = 8'b10011100;
DRAM[5624] = 8'b10011100;
DRAM[5625] = 8'b10011011;
DRAM[5626] = 8'b10011010;
DRAM[5627] = 8'b10011011;
DRAM[5628] = 8'b10011100;
DRAM[5629] = 8'b10011101;
DRAM[5630] = 8'b10011001;
DRAM[5631] = 8'b10011001;
DRAM[5632] = 8'b01100010;
DRAM[5633] = 8'b01100010;
DRAM[5634] = 8'b01100010;
DRAM[5635] = 8'b01100010;
DRAM[5636] = 8'b01100100;
DRAM[5637] = 8'b01101011;
DRAM[5638] = 8'b01111000;
DRAM[5639] = 8'b10001111;
DRAM[5640] = 8'b10011111;
DRAM[5641] = 8'b10101001;
DRAM[5642] = 8'b10101100;
DRAM[5643] = 8'b10101111;
DRAM[5644] = 8'b10101110;
DRAM[5645] = 8'b10100110;
DRAM[5646] = 8'b10010011;
DRAM[5647] = 8'b01101111;
DRAM[5648] = 8'b01001110;
DRAM[5649] = 8'b01001101;
DRAM[5650] = 8'b01010110;
DRAM[5651] = 8'b01011110;
DRAM[5652] = 8'b01100010;
DRAM[5653] = 8'b01100011;
DRAM[5654] = 8'b01100010;
DRAM[5655] = 8'b01100101;
DRAM[5656] = 8'b01100010;
DRAM[5657] = 8'b01100100;
DRAM[5658] = 8'b01100010;
DRAM[5659] = 8'b01011100;
DRAM[5660] = 8'b01010100;
DRAM[5661] = 8'b10011011;
DRAM[5662] = 8'b11001110;
DRAM[5663] = 8'b11000010;
DRAM[5664] = 8'b10111000;
DRAM[5665] = 8'b10100100;
DRAM[5666] = 8'b10000110;
DRAM[5667] = 8'b10011001;
DRAM[5668] = 8'b10010011;
DRAM[5669] = 8'b01110001;
DRAM[5670] = 8'b01111001;
DRAM[5671] = 8'b01111010;
DRAM[5672] = 8'b01110001;
DRAM[5673] = 8'b01110100;
DRAM[5674] = 8'b10001001;
DRAM[5675] = 8'b10001011;
DRAM[5676] = 8'b10000111;
DRAM[5677] = 8'b01111100;
DRAM[5678] = 8'b01111100;
DRAM[5679] = 8'b10000001;
DRAM[5680] = 8'b10000101;
DRAM[5681] = 8'b10000100;
DRAM[5682] = 8'b10001101;
DRAM[5683] = 8'b10001101;
DRAM[5684] = 8'b10001001;
DRAM[5685] = 8'b10000001;
DRAM[5686] = 8'b10001100;
DRAM[5687] = 8'b01101110;
DRAM[5688] = 8'b01101100;
DRAM[5689] = 8'b01010110;
DRAM[5690] = 8'b01010000;
DRAM[5691] = 8'b01100010;
DRAM[5692] = 8'b10011100;
DRAM[5693] = 8'b10011001;
DRAM[5694] = 8'b01111110;
DRAM[5695] = 8'b01110000;
DRAM[5696] = 8'b01100110;
DRAM[5697] = 8'b01010000;
DRAM[5698] = 8'b01011011;
DRAM[5699] = 8'b01010000;
DRAM[5700] = 8'b01001100;
DRAM[5701] = 8'b00111111;
DRAM[5702] = 8'b00110100;
DRAM[5703] = 8'b00111011;
DRAM[5704] = 8'b00110100;
DRAM[5705] = 8'b10110110;
DRAM[5706] = 8'b10100100;
DRAM[5707] = 8'b10100101;
DRAM[5708] = 8'b11000000;
DRAM[5709] = 8'b11000010;
DRAM[5710] = 8'b11000101;
DRAM[5711] = 8'b11000000;
DRAM[5712] = 8'b11000100;
DRAM[5713] = 8'b11000100;
DRAM[5714] = 8'b11000000;
DRAM[5715] = 8'b11000010;
DRAM[5716] = 8'b11000101;
DRAM[5717] = 8'b11001001;
DRAM[5718] = 8'b11000111;
DRAM[5719] = 8'b11001001;
DRAM[5720] = 8'b11001010;
DRAM[5721] = 8'b11001100;
DRAM[5722] = 8'b11001011;
DRAM[5723] = 8'b11001100;
DRAM[5724] = 8'b11010000;
DRAM[5725] = 8'b10110010;
DRAM[5726] = 8'b01111111;
DRAM[5727] = 8'b01011001;
DRAM[5728] = 8'b01010110;
DRAM[5729] = 8'b01011111;
DRAM[5730] = 8'b10000101;
DRAM[5731] = 8'b11000110;
DRAM[5732] = 8'b10110100;
DRAM[5733] = 8'b00100010;
DRAM[5734] = 8'b00101010;
DRAM[5735] = 8'b00110011;
DRAM[5736] = 8'b00110001;
DRAM[5737] = 8'b00101100;
DRAM[5738] = 8'b00110000;
DRAM[5739] = 8'b00110001;
DRAM[5740] = 8'b00101111;
DRAM[5741] = 8'b01101000;
DRAM[5742] = 8'b10010111;
DRAM[5743] = 8'b10010001;
DRAM[5744] = 8'b10010110;
DRAM[5745] = 8'b10100000;
DRAM[5746] = 8'b10100000;
DRAM[5747] = 8'b10011111;
DRAM[5748] = 8'b10011110;
DRAM[5749] = 8'b10011110;
DRAM[5750] = 8'b10011011;
DRAM[5751] = 8'b10011011;
DRAM[5752] = 8'b10011100;
DRAM[5753] = 8'b10011011;
DRAM[5754] = 8'b10011010;
DRAM[5755] = 8'b10011001;
DRAM[5756] = 8'b10011001;
DRAM[5757] = 8'b10011010;
DRAM[5758] = 8'b10011001;
DRAM[5759] = 8'b10011001;
DRAM[5760] = 8'b01100010;
DRAM[5761] = 8'b01101000;
DRAM[5762] = 8'b01100011;
DRAM[5763] = 8'b01100010;
DRAM[5764] = 8'b01100110;
DRAM[5765] = 8'b01101110;
DRAM[5766] = 8'b01111000;
DRAM[5767] = 8'b10010000;
DRAM[5768] = 8'b10011111;
DRAM[5769] = 8'b10101100;
DRAM[5770] = 8'b10101011;
DRAM[5771] = 8'b10101101;
DRAM[5772] = 8'b10101110;
DRAM[5773] = 8'b10100111;
DRAM[5774] = 8'b10010011;
DRAM[5775] = 8'b01110000;
DRAM[5776] = 8'b01001110;
DRAM[5777] = 8'b01001110;
DRAM[5778] = 8'b01011000;
DRAM[5779] = 8'b01011111;
DRAM[5780] = 8'b01011111;
DRAM[5781] = 8'b01100011;
DRAM[5782] = 8'b01100000;
DRAM[5783] = 8'b01101001;
DRAM[5784] = 8'b01100010;
DRAM[5785] = 8'b01100010;
DRAM[5786] = 8'b01100101;
DRAM[5787] = 8'b01100001;
DRAM[5788] = 8'b01011011;
DRAM[5789] = 8'b01110101;
DRAM[5790] = 8'b11010000;
DRAM[5791] = 8'b11000110;
DRAM[5792] = 8'b11000011;
DRAM[5793] = 8'b10011110;
DRAM[5794] = 8'b01111100;
DRAM[5795] = 8'b10000011;
DRAM[5796] = 8'b01110110;
DRAM[5797] = 8'b01110001;
DRAM[5798] = 8'b01110110;
DRAM[5799] = 8'b01110010;
DRAM[5800] = 8'b01110000;
DRAM[5801] = 8'b10000111;
DRAM[5802] = 8'b10001000;
DRAM[5803] = 8'b10000110;
DRAM[5804] = 8'b01111001;
DRAM[5805] = 8'b10000011;
DRAM[5806] = 8'b10000101;
DRAM[5807] = 8'b10000110;
DRAM[5808] = 8'b10000011;
DRAM[5809] = 8'b10001000;
DRAM[5810] = 8'b10001101;
DRAM[5811] = 8'b10000101;
DRAM[5812] = 8'b01110101;
DRAM[5813] = 8'b10001010;
DRAM[5814] = 8'b01110111;
DRAM[5815] = 8'b01110110;
DRAM[5816] = 8'b01100111;
DRAM[5817] = 8'b01111100;
DRAM[5818] = 8'b01100010;
DRAM[5819] = 8'b01101001;
DRAM[5820] = 8'b01100000;
DRAM[5821] = 8'b01111010;
DRAM[5822] = 8'b01011010;
DRAM[5823] = 8'b00111110;
DRAM[5824] = 8'b01001111;
DRAM[5825] = 8'b01010110;
DRAM[5826] = 8'b01000010;
DRAM[5827] = 8'b01001000;
DRAM[5828] = 8'b00101100;
DRAM[5829] = 8'b00100111;
DRAM[5830] = 8'b00101000;
DRAM[5831] = 8'b01000110;
DRAM[5832] = 8'b10011011;
DRAM[5833] = 8'b10011110;
DRAM[5834] = 8'b10110100;
DRAM[5835] = 8'b11001010;
DRAM[5836] = 8'b11000111;
DRAM[5837] = 8'b11000010;
DRAM[5838] = 8'b11000001;
DRAM[5839] = 8'b11000001;
DRAM[5840] = 8'b11000100;
DRAM[5841] = 8'b11000001;
DRAM[5842] = 8'b10111111;
DRAM[5843] = 8'b11000100;
DRAM[5844] = 8'b11000110;
DRAM[5845] = 8'b11000111;
DRAM[5846] = 8'b11001000;
DRAM[5847] = 8'b11000101;
DRAM[5848] = 8'b11001110;
DRAM[5849] = 8'b11001101;
DRAM[5850] = 8'b11001100;
DRAM[5851] = 8'b10010111;
DRAM[5852] = 8'b01101100;
DRAM[5853] = 8'b01011001;
DRAM[5854] = 8'b01011110;
DRAM[5855] = 8'b01011001;
DRAM[5856] = 8'b01101000;
DRAM[5857] = 8'b10000111;
DRAM[5858] = 8'b10111010;
DRAM[5859] = 8'b11001010;
DRAM[5860] = 8'b01001001;
DRAM[5861] = 8'b00100110;
DRAM[5862] = 8'b00110010;
DRAM[5863] = 8'b00110011;
DRAM[5864] = 8'b00110100;
DRAM[5865] = 8'b00101110;
DRAM[5866] = 8'b00111001;
DRAM[5867] = 8'b00101100;
DRAM[5868] = 8'b00111001;
DRAM[5869] = 8'b10001010;
DRAM[5870] = 8'b10010010;
DRAM[5871] = 8'b10010000;
DRAM[5872] = 8'b10011110;
DRAM[5873] = 8'b10100001;
DRAM[5874] = 8'b10100001;
DRAM[5875] = 8'b10100001;
DRAM[5876] = 8'b10011110;
DRAM[5877] = 8'b10011111;
DRAM[5878] = 8'b10011111;
DRAM[5879] = 8'b10011101;
DRAM[5880] = 8'b10011011;
DRAM[5881] = 8'b10011001;
DRAM[5882] = 8'b10011011;
DRAM[5883] = 8'b10011011;
DRAM[5884] = 8'b10011001;
DRAM[5885] = 8'b10011001;
DRAM[5886] = 8'b10011000;
DRAM[5887] = 8'b10011011;
DRAM[5888] = 8'b01100110;
DRAM[5889] = 8'b01100101;
DRAM[5890] = 8'b01100100;
DRAM[5891] = 8'b01011110;
DRAM[5892] = 8'b01101000;
DRAM[5893] = 8'b01101100;
DRAM[5894] = 8'b01111011;
DRAM[5895] = 8'b10001101;
DRAM[5896] = 8'b10100000;
DRAM[5897] = 8'b10101011;
DRAM[5898] = 8'b10101100;
DRAM[5899] = 8'b10101110;
DRAM[5900] = 8'b10101100;
DRAM[5901] = 8'b10100110;
DRAM[5902] = 8'b10010011;
DRAM[5903] = 8'b01101110;
DRAM[5904] = 8'b01001100;
DRAM[5905] = 8'b01001101;
DRAM[5906] = 8'b01011001;
DRAM[5907] = 8'b01100010;
DRAM[5908] = 8'b01100010;
DRAM[5909] = 8'b01100011;
DRAM[5910] = 8'b01100010;
DRAM[5911] = 8'b01100101;
DRAM[5912] = 8'b01100010;
DRAM[5913] = 8'b01100101;
DRAM[5914] = 8'b01100000;
DRAM[5915] = 8'b01100000;
DRAM[5916] = 8'b01011000;
DRAM[5917] = 8'b01001110;
DRAM[5918] = 8'b11011000;
DRAM[5919] = 8'b11001010;
DRAM[5920] = 8'b11000110;
DRAM[5921] = 8'b10100010;
DRAM[5922] = 8'b01110111;
DRAM[5923] = 8'b10001101;
DRAM[5924] = 8'b10001011;
DRAM[5925] = 8'b01111011;
DRAM[5926] = 8'b01110000;
DRAM[5927] = 8'b01101101;
DRAM[5928] = 8'b10000000;
DRAM[5929] = 8'b10001000;
DRAM[5930] = 8'b10001001;
DRAM[5931] = 8'b01111011;
DRAM[5932] = 8'b01111111;
DRAM[5933] = 8'b10000100;
DRAM[5934] = 8'b10000101;
DRAM[5935] = 8'b10000001;
DRAM[5936] = 8'b10000010;
DRAM[5937] = 8'b10001110;
DRAM[5938] = 8'b10000011;
DRAM[5939] = 8'b01110100;
DRAM[5940] = 8'b10000110;
DRAM[5941] = 8'b01110111;
DRAM[5942] = 8'b01110011;
DRAM[5943] = 8'b01110101;
DRAM[5944] = 8'b01011011;
DRAM[5945] = 8'b00111101;
DRAM[5946] = 8'b00111001;
DRAM[5947] = 8'b00111001;
DRAM[5948] = 8'b01011011;
DRAM[5949] = 8'b01110000;
DRAM[5950] = 8'b01011110;
DRAM[5951] = 8'b01100011;
DRAM[5952] = 8'b01100011;
DRAM[5953] = 8'b01000100;
DRAM[5954] = 8'b00111000;
DRAM[5955] = 8'b01000011;
DRAM[5956] = 8'b00100111;
DRAM[5957] = 8'b00100110;
DRAM[5958] = 8'b01000100;
DRAM[5959] = 8'b10100001;
DRAM[5960] = 8'b10001000;
DRAM[5961] = 8'b10110111;
DRAM[5962] = 8'b10111010;
DRAM[5963] = 8'b11000001;
DRAM[5964] = 8'b11000100;
DRAM[5965] = 8'b11000001;
DRAM[5966] = 8'b11000010;
DRAM[5967] = 8'b10111110;
DRAM[5968] = 8'b11000010;
DRAM[5969] = 8'b11000000;
DRAM[5970] = 8'b10111110;
DRAM[5971] = 8'b11000000;
DRAM[5972] = 8'b11000100;
DRAM[5973] = 8'b11000101;
DRAM[5974] = 8'b11001010;
DRAM[5975] = 8'b11001010;
DRAM[5976] = 8'b11001111;
DRAM[5977] = 8'b10100110;
DRAM[5978] = 8'b01010110;
DRAM[5979] = 8'b01011101;
DRAM[5980] = 8'b01011000;
DRAM[5981] = 8'b01011010;
DRAM[5982] = 8'b01101000;
DRAM[5983] = 8'b01111110;
DRAM[5984] = 8'b10100011;
DRAM[5985] = 8'b11000000;
DRAM[5986] = 8'b10100101;
DRAM[5987] = 8'b00101000;
DRAM[5988] = 8'b00101010;
DRAM[5989] = 8'b00101110;
DRAM[5990] = 8'b00110011;
DRAM[5991] = 8'b00101110;
DRAM[5992] = 8'b00101100;
DRAM[5993] = 8'b00110000;
DRAM[5994] = 8'b00110101;
DRAM[5995] = 8'b00101101;
DRAM[5996] = 8'b01011101;
DRAM[5997] = 8'b10010011;
DRAM[5998] = 8'b10010001;
DRAM[5999] = 8'b10011000;
DRAM[6000] = 8'b10100001;
DRAM[6001] = 8'b10100100;
DRAM[6002] = 8'b10100001;
DRAM[6003] = 8'b10100000;
DRAM[6004] = 8'b10011110;
DRAM[6005] = 8'b10011110;
DRAM[6006] = 8'b10011110;
DRAM[6007] = 8'b10011101;
DRAM[6008] = 8'b10011100;
DRAM[6009] = 8'b10011011;
DRAM[6010] = 8'b10011001;
DRAM[6011] = 8'b10011001;
DRAM[6012] = 8'b10011100;
DRAM[6013] = 8'b10011000;
DRAM[6014] = 8'b10011001;
DRAM[6015] = 8'b10011010;
DRAM[6016] = 8'b01101001;
DRAM[6017] = 8'b01101001;
DRAM[6018] = 8'b01100100;
DRAM[6019] = 8'b01100011;
DRAM[6020] = 8'b01100101;
DRAM[6021] = 8'b01101010;
DRAM[6022] = 8'b01110111;
DRAM[6023] = 8'b10001101;
DRAM[6024] = 8'b10011011;
DRAM[6025] = 8'b10101001;
DRAM[6026] = 8'b10101100;
DRAM[6027] = 8'b10101010;
DRAM[6028] = 8'b10101011;
DRAM[6029] = 8'b10100101;
DRAM[6030] = 8'b10010101;
DRAM[6031] = 8'b01101111;
DRAM[6032] = 8'b01010000;
DRAM[6033] = 8'b01001100;
DRAM[6034] = 8'b01010111;
DRAM[6035] = 8'b01011111;
DRAM[6036] = 8'b01100001;
DRAM[6037] = 8'b01100000;
DRAM[6038] = 8'b01100011;
DRAM[6039] = 8'b01100100;
DRAM[6040] = 8'b01100010;
DRAM[6041] = 8'b01100100;
DRAM[6042] = 8'b01100100;
DRAM[6043] = 8'b01100001;
DRAM[6044] = 8'b01011110;
DRAM[6045] = 8'b01010000;
DRAM[6046] = 8'b10111111;
DRAM[6047] = 8'b11001001;
DRAM[6048] = 8'b11000110;
DRAM[6049] = 8'b10100110;
DRAM[6050] = 8'b10000100;
DRAM[6051] = 8'b10001100;
DRAM[6052] = 8'b10011001;
DRAM[6053] = 8'b01111110;
DRAM[6054] = 8'b01101011;
DRAM[6055] = 8'b01110111;
DRAM[6056] = 8'b10000111;
DRAM[6057] = 8'b10000111;
DRAM[6058] = 8'b01111010;
DRAM[6059] = 8'b01111100;
DRAM[6060] = 8'b01111101;
DRAM[6061] = 8'b10001000;
DRAM[6062] = 8'b01111111;
DRAM[6063] = 8'b10000010;
DRAM[6064] = 8'b10001011;
DRAM[6065] = 8'b10001000;
DRAM[6066] = 8'b01101000;
DRAM[6067] = 8'b10000101;
DRAM[6068] = 8'b01111111;
DRAM[6069] = 8'b01100111;
DRAM[6070] = 8'b01000110;
DRAM[6071] = 8'b01010100;
DRAM[6072] = 8'b01000101;
DRAM[6073] = 8'b00111000;
DRAM[6074] = 8'b00110101;
DRAM[6075] = 8'b01010110;
DRAM[6076] = 8'b01101110;
DRAM[6077] = 8'b01011000;
DRAM[6078] = 8'b00110000;
DRAM[6079] = 8'b01100011;
DRAM[6080] = 8'b01011100;
DRAM[6081] = 8'b01010010;
DRAM[6082] = 8'b00110111;
DRAM[6083] = 8'b01010010;
DRAM[6084] = 8'b00011111;
DRAM[6085] = 8'b01100001;
DRAM[6086] = 8'b10100000;
DRAM[6087] = 8'b10000100;
DRAM[6088] = 8'b10110110;
DRAM[6089] = 8'b10111110;
DRAM[6090] = 8'b10110010;
DRAM[6091] = 8'b10111010;
DRAM[6092] = 8'b10111111;
DRAM[6093] = 8'b10111111;
DRAM[6094] = 8'b10111101;
DRAM[6095] = 8'b10111010;
DRAM[6096] = 8'b10111110;
DRAM[6097] = 8'b10111110;
DRAM[6098] = 8'b11000001;
DRAM[6099] = 8'b11000010;
DRAM[6100] = 8'b11000100;
DRAM[6101] = 8'b11000101;
DRAM[6102] = 8'b11000111;
DRAM[6103] = 8'b10100111;
DRAM[6104] = 8'b01110101;
DRAM[6105] = 8'b10000011;
DRAM[6106] = 8'b01100010;
DRAM[6107] = 8'b01100000;
DRAM[6108] = 8'b01101110;
DRAM[6109] = 8'b10000110;
DRAM[6110] = 8'b10011101;
DRAM[6111] = 8'b10101010;
DRAM[6112] = 8'b10111001;
DRAM[6113] = 8'b10101110;
DRAM[6114] = 8'b00110100;
DRAM[6115] = 8'b00110010;
DRAM[6116] = 8'b00110011;
DRAM[6117] = 8'b00110110;
DRAM[6118] = 8'b00110011;
DRAM[6119] = 8'b00101100;
DRAM[6120] = 8'b00101101;
DRAM[6121] = 8'b01000000;
DRAM[6122] = 8'b00111000;
DRAM[6123] = 8'b00111100;
DRAM[6124] = 8'b10000100;
DRAM[6125] = 8'b10010101;
DRAM[6126] = 8'b10010000;
DRAM[6127] = 8'b10100000;
DRAM[6128] = 8'b10100101;
DRAM[6129] = 8'b10100011;
DRAM[6130] = 8'b10100001;
DRAM[6131] = 8'b10100010;
DRAM[6132] = 8'b10100010;
DRAM[6133] = 8'b10011110;
DRAM[6134] = 8'b10011110;
DRAM[6135] = 8'b10011101;
DRAM[6136] = 8'b10011100;
DRAM[6137] = 8'b10011011;
DRAM[6138] = 8'b10011101;
DRAM[6139] = 8'b10011100;
DRAM[6140] = 8'b10011010;
DRAM[6141] = 8'b10011011;
DRAM[6142] = 8'b10011010;
DRAM[6143] = 8'b10011001;
DRAM[6144] = 8'b01101001;
DRAM[6145] = 8'b01101010;
DRAM[6146] = 8'b01100111;
DRAM[6147] = 8'b01100011;
DRAM[6148] = 8'b01100011;
DRAM[6149] = 8'b01101000;
DRAM[6150] = 8'b01110110;
DRAM[6151] = 8'b10001100;
DRAM[6152] = 8'b10011110;
DRAM[6153] = 8'b10101010;
DRAM[6154] = 8'b10101100;
DRAM[6155] = 8'b10101100;
DRAM[6156] = 8'b10101010;
DRAM[6157] = 8'b10100111;
DRAM[6158] = 8'b10010011;
DRAM[6159] = 8'b01110100;
DRAM[6160] = 8'b01001110;
DRAM[6161] = 8'b01001110;
DRAM[6162] = 8'b01010111;
DRAM[6163] = 8'b01100000;
DRAM[6164] = 8'b01100000;
DRAM[6165] = 8'b01100000;
DRAM[6166] = 8'b01100011;
DRAM[6167] = 8'b01100100;
DRAM[6168] = 8'b01100100;
DRAM[6169] = 8'b01100100;
DRAM[6170] = 8'b01100000;
DRAM[6171] = 8'b01100101;
DRAM[6172] = 8'b01100010;
DRAM[6173] = 8'b01010100;
DRAM[6174] = 8'b10011100;
DRAM[6175] = 8'b11001010;
DRAM[6176] = 8'b11000010;
DRAM[6177] = 8'b10111000;
DRAM[6178] = 8'b10011100;
DRAM[6179] = 8'b10001011;
DRAM[6180] = 8'b10001000;
DRAM[6181] = 8'b01101101;
DRAM[6182] = 8'b01110100;
DRAM[6183] = 8'b10001001;
DRAM[6184] = 8'b10000110;
DRAM[6185] = 8'b01110111;
DRAM[6186] = 8'b01110111;
DRAM[6187] = 8'b10000000;
DRAM[6188] = 8'b10000000;
DRAM[6189] = 8'b01111111;
DRAM[6190] = 8'b01110101;
DRAM[6191] = 8'b10001001;
DRAM[6192] = 8'b10001000;
DRAM[6193] = 8'b10001110;
DRAM[6194] = 8'b01101100;
DRAM[6195] = 8'b01111100;
DRAM[6196] = 8'b01001010;
DRAM[6197] = 8'b01000100;
DRAM[6198] = 8'b01010000;
DRAM[6199] = 8'b00110111;
DRAM[6200] = 8'b00110100;
DRAM[6201] = 8'b00110000;
DRAM[6202] = 8'b00110001;
DRAM[6203] = 8'b01110001;
DRAM[6204] = 8'b01011010;
DRAM[6205] = 8'b00110001;
DRAM[6206] = 8'b01001010;
DRAM[6207] = 8'b01010101;
DRAM[6208] = 8'b01011010;
DRAM[6209] = 8'b00110011;
DRAM[6210] = 8'b00100101;
DRAM[6211] = 8'b01011111;
DRAM[6212] = 8'b01110100;
DRAM[6213] = 8'b10010010;
DRAM[6214] = 8'b10001110;
DRAM[6215] = 8'b11000010;
DRAM[6216] = 8'b10111101;
DRAM[6217] = 8'b10110101;
DRAM[6218] = 8'b10110101;
DRAM[6219] = 8'b10111010;
DRAM[6220] = 8'b10111001;
DRAM[6221] = 8'b10111001;
DRAM[6222] = 8'b10110111;
DRAM[6223] = 8'b10111011;
DRAM[6224] = 8'b10111101;
DRAM[6225] = 8'b10111111;
DRAM[6226] = 8'b11000001;
DRAM[6227] = 8'b11000011;
DRAM[6228] = 8'b11000110;
DRAM[6229] = 8'b10101011;
DRAM[6230] = 8'b01101100;
DRAM[6231] = 8'b01011010;
DRAM[6232] = 8'b01101010;
DRAM[6233] = 8'b10001101;
DRAM[6234] = 8'b10010100;
DRAM[6235] = 8'b10011101;
DRAM[6236] = 8'b10100101;
DRAM[6237] = 8'b10100110;
DRAM[6238] = 8'b10101010;
DRAM[6239] = 8'b10110101;
DRAM[6240] = 8'b10110111;
DRAM[6241] = 8'b00101101;
DRAM[6242] = 8'b00101011;
DRAM[6243] = 8'b00110011;
DRAM[6244] = 8'b00111000;
DRAM[6245] = 8'b00110010;
DRAM[6246] = 8'b00110010;
DRAM[6247] = 8'b00110100;
DRAM[6248] = 8'b00101100;
DRAM[6249] = 8'b00110111;
DRAM[6250] = 8'b00110000;
DRAM[6251] = 8'b01010101;
DRAM[6252] = 8'b10010000;
DRAM[6253] = 8'b10010010;
DRAM[6254] = 8'b10010101;
DRAM[6255] = 8'b10100101;
DRAM[6256] = 8'b10100011;
DRAM[6257] = 8'b10100100;
DRAM[6258] = 8'b10100100;
DRAM[6259] = 8'b10100011;
DRAM[6260] = 8'b10100010;
DRAM[6261] = 8'b10100000;
DRAM[6262] = 8'b10011101;
DRAM[6263] = 8'b10011101;
DRAM[6264] = 8'b10011101;
DRAM[6265] = 8'b10011001;
DRAM[6266] = 8'b10011010;
DRAM[6267] = 8'b10011011;
DRAM[6268] = 8'b10011010;
DRAM[6269] = 8'b10011100;
DRAM[6270] = 8'b10011000;
DRAM[6271] = 8'b10010111;
DRAM[6272] = 8'b01101100;
DRAM[6273] = 8'b01101000;
DRAM[6274] = 8'b01100101;
DRAM[6275] = 8'b01101000;
DRAM[6276] = 8'b01100110;
DRAM[6277] = 8'b01100111;
DRAM[6278] = 8'b01110110;
DRAM[6279] = 8'b10001101;
DRAM[6280] = 8'b10011110;
DRAM[6281] = 8'b10101010;
DRAM[6282] = 8'b10101011;
DRAM[6283] = 8'b10101101;
DRAM[6284] = 8'b10101100;
DRAM[6285] = 8'b10100110;
DRAM[6286] = 8'b10010100;
DRAM[6287] = 8'b01110110;
DRAM[6288] = 8'b01001110;
DRAM[6289] = 8'b01001110;
DRAM[6290] = 8'b01011001;
DRAM[6291] = 8'b01011100;
DRAM[6292] = 8'b01100001;
DRAM[6293] = 8'b01100000;
DRAM[6294] = 8'b01100010;
DRAM[6295] = 8'b01100011;
DRAM[6296] = 8'b01100000;
DRAM[6297] = 8'b01100101;
DRAM[6298] = 8'b01100001;
DRAM[6299] = 8'b01100110;
DRAM[6300] = 8'b01100110;
DRAM[6301] = 8'b01011100;
DRAM[6302] = 8'b01101110;
DRAM[6303] = 8'b11010101;
DRAM[6304] = 8'b11000111;
DRAM[6305] = 8'b11000010;
DRAM[6306] = 8'b10100111;
DRAM[6307] = 8'b10011111;
DRAM[6308] = 8'b01111101;
DRAM[6309] = 8'b01110010;
DRAM[6310] = 8'b10000001;
DRAM[6311] = 8'b10001000;
DRAM[6312] = 8'b01111110;
DRAM[6313] = 8'b01110011;
DRAM[6314] = 8'b01111100;
DRAM[6315] = 8'b01111110;
DRAM[6316] = 8'b01111101;
DRAM[6317] = 8'b01111000;
DRAM[6318] = 8'b10001000;
DRAM[6319] = 8'b01111111;
DRAM[6320] = 8'b01100100;
DRAM[6321] = 8'b01101100;
DRAM[6322] = 8'b01100111;
DRAM[6323] = 8'b01000010;
DRAM[6324] = 8'b01001010;
DRAM[6325] = 8'b01001001;
DRAM[6326] = 8'b00111011;
DRAM[6327] = 8'b00111000;
DRAM[6328] = 8'b00110100;
DRAM[6329] = 8'b00101100;
DRAM[6330] = 8'b01010101;
DRAM[6331] = 8'b01001010;
DRAM[6332] = 8'b00111011;
DRAM[6333] = 8'b01000111;
DRAM[6334] = 8'b01100110;
DRAM[6335] = 8'b01101011;
DRAM[6336] = 8'b00110001;
DRAM[6337] = 8'b01000011;
DRAM[6338] = 8'b00111101;
DRAM[6339] = 8'b10000010;
DRAM[6340] = 8'b10001100;
DRAM[6341] = 8'b10010011;
DRAM[6342] = 8'b11000000;
DRAM[6343] = 8'b11000011;
DRAM[6344] = 8'b10110100;
DRAM[6345] = 8'b10110011;
DRAM[6346] = 8'b10110101;
DRAM[6347] = 8'b10110111;
DRAM[6348] = 8'b10110011;
DRAM[6349] = 8'b10110010;
DRAM[6350] = 8'b10110100;
DRAM[6351] = 8'b10111011;
DRAM[6352] = 8'b10111110;
DRAM[6353] = 8'b10111111;
DRAM[6354] = 8'b11000001;
DRAM[6355] = 8'b11000101;
DRAM[6356] = 8'b01100010;
DRAM[6357] = 8'b01010100;
DRAM[6358] = 8'b01001100;
DRAM[6359] = 8'b01111011;
DRAM[6360] = 8'b01110000;
DRAM[6361] = 8'b10000010;
DRAM[6362] = 8'b10100010;
DRAM[6363] = 8'b10100111;
DRAM[6364] = 8'b10101000;
DRAM[6365] = 8'b10101101;
DRAM[6366] = 8'b10111010;
DRAM[6367] = 8'b11000000;
DRAM[6368] = 8'b00111000;
DRAM[6369] = 8'b00101001;
DRAM[6370] = 8'b00101111;
DRAM[6371] = 8'b00110101;
DRAM[6372] = 8'b00110111;
DRAM[6373] = 8'b00110110;
DRAM[6374] = 8'b00110001;
DRAM[6375] = 8'b00101110;
DRAM[6376] = 8'b00110101;
DRAM[6377] = 8'b00110110;
DRAM[6378] = 8'b00110100;
DRAM[6379] = 8'b01110010;
DRAM[6380] = 8'b10010011;
DRAM[6381] = 8'b10001110;
DRAM[6382] = 8'b10011110;
DRAM[6383] = 8'b10100101;
DRAM[6384] = 8'b10100110;
DRAM[6385] = 8'b10100101;
DRAM[6386] = 8'b10100100;
DRAM[6387] = 8'b10100100;
DRAM[6388] = 8'b10100001;
DRAM[6389] = 8'b10011111;
DRAM[6390] = 8'b10011111;
DRAM[6391] = 8'b10011110;
DRAM[6392] = 8'b10011011;
DRAM[6393] = 8'b10011100;
DRAM[6394] = 8'b10011011;
DRAM[6395] = 8'b10011101;
DRAM[6396] = 8'b10011011;
DRAM[6397] = 8'b10011000;
DRAM[6398] = 8'b10011010;
DRAM[6399] = 8'b10010111;
DRAM[6400] = 8'b01101110;
DRAM[6401] = 8'b01101000;
DRAM[6402] = 8'b01100111;
DRAM[6403] = 8'b01100100;
DRAM[6404] = 8'b01100011;
DRAM[6405] = 8'b01100111;
DRAM[6406] = 8'b01110011;
DRAM[6407] = 8'b10001000;
DRAM[6408] = 8'b10011111;
DRAM[6409] = 8'b10101010;
DRAM[6410] = 8'b10101010;
DRAM[6411] = 8'b10101110;
DRAM[6412] = 8'b10101011;
DRAM[6413] = 8'b10100110;
DRAM[6414] = 8'b10010101;
DRAM[6415] = 8'b01110101;
DRAM[6416] = 8'b01001100;
DRAM[6417] = 8'b01001011;
DRAM[6418] = 8'b01011000;
DRAM[6419] = 8'b01011100;
DRAM[6420] = 8'b01100001;
DRAM[6421] = 8'b01011111;
DRAM[6422] = 8'b01100010;
DRAM[6423] = 8'b01100000;
DRAM[6424] = 8'b01100001;
DRAM[6425] = 8'b01100010;
DRAM[6426] = 8'b01100010;
DRAM[6427] = 8'b01100111;
DRAM[6428] = 8'b01101000;
DRAM[6429] = 8'b01100101;
DRAM[6430] = 8'b01010110;
DRAM[6431] = 8'b10101101;
DRAM[6432] = 8'b11010001;
DRAM[6433] = 8'b10111110;
DRAM[6434] = 8'b10100111;
DRAM[6435] = 8'b10110000;
DRAM[6436] = 8'b01100010;
DRAM[6437] = 8'b10000100;
DRAM[6438] = 8'b10000000;
DRAM[6439] = 8'b01111100;
DRAM[6440] = 8'b01101110;
DRAM[6441] = 8'b10000001;
DRAM[6442] = 8'b01111101;
DRAM[6443] = 8'b01111000;
DRAM[6444] = 8'b01111010;
DRAM[6445] = 8'b10000100;
DRAM[6446] = 8'b01111110;
DRAM[6447] = 8'b01110100;
DRAM[6448] = 8'b01001010;
DRAM[6449] = 8'b01001010;
DRAM[6450] = 8'b01001100;
DRAM[6451] = 8'b01001011;
DRAM[6452] = 8'b01001101;
DRAM[6453] = 8'b00111010;
DRAM[6454] = 8'b00110000;
DRAM[6455] = 8'b01011111;
DRAM[6456] = 8'b00101000;
DRAM[6457] = 8'b00111101;
DRAM[6458] = 8'b01100111;
DRAM[6459] = 8'b00101001;
DRAM[6460] = 8'b00111000;
DRAM[6461] = 8'b00111101;
DRAM[6462] = 8'b01000111;
DRAM[6463] = 8'b01001010;
DRAM[6464] = 8'b01011110;
DRAM[6465] = 8'b00111011;
DRAM[6466] = 8'b01110010;
DRAM[6467] = 8'b01111110;
DRAM[6468] = 8'b10010111;
DRAM[6469] = 8'b11000011;
DRAM[6470] = 8'b11000010;
DRAM[6471] = 8'b10111110;
DRAM[6472] = 8'b10110110;
DRAM[6473] = 8'b10110100;
DRAM[6474] = 8'b10110101;
DRAM[6475] = 8'b10110100;
DRAM[6476] = 8'b10101100;
DRAM[6477] = 8'b10110011;
DRAM[6478] = 8'b10110001;
DRAM[6479] = 8'b10111101;
DRAM[6480] = 8'b10111111;
DRAM[6481] = 8'b10111101;
DRAM[6482] = 8'b10111001;
DRAM[6483] = 8'b10000010;
DRAM[6484] = 8'b01001001;
DRAM[6485] = 8'b01010001;
DRAM[6486] = 8'b01100101;
DRAM[6487] = 8'b01110111;
DRAM[6488] = 8'b01111010;
DRAM[6489] = 8'b01110000;
DRAM[6490] = 8'b10011000;
DRAM[6491] = 8'b10100111;
DRAM[6492] = 8'b10101101;
DRAM[6493] = 8'b11000000;
DRAM[6494] = 8'b10011000;
DRAM[6495] = 8'b00100100;
DRAM[6496] = 8'b00101110;
DRAM[6497] = 8'b00101101;
DRAM[6498] = 8'b00110000;
DRAM[6499] = 8'b00110101;
DRAM[6500] = 8'b00111010;
DRAM[6501] = 8'b00110110;
DRAM[6502] = 8'b00101111;
DRAM[6503] = 8'b00101010;
DRAM[6504] = 8'b00110011;
DRAM[6505] = 8'b00110001;
DRAM[6506] = 8'b01001001;
DRAM[6507] = 8'b10000100;
DRAM[6508] = 8'b10001011;
DRAM[6509] = 8'b10001111;
DRAM[6510] = 8'b10100101;
DRAM[6511] = 8'b10101000;
DRAM[6512] = 8'b10100100;
DRAM[6513] = 8'b10100101;
DRAM[6514] = 8'b10100000;
DRAM[6515] = 8'b10100101;
DRAM[6516] = 8'b10100010;
DRAM[6517] = 8'b10100001;
DRAM[6518] = 8'b10100000;
DRAM[6519] = 8'b10011110;
DRAM[6520] = 8'b10011101;
DRAM[6521] = 8'b10011110;
DRAM[6522] = 8'b10011110;
DRAM[6523] = 8'b10011100;
DRAM[6524] = 8'b10011100;
DRAM[6525] = 8'b10011000;
DRAM[6526] = 8'b10011000;
DRAM[6527] = 8'b10010111;
DRAM[6528] = 8'b01101011;
DRAM[6529] = 8'b01101101;
DRAM[6530] = 8'b01100110;
DRAM[6531] = 8'b01100101;
DRAM[6532] = 8'b01100011;
DRAM[6533] = 8'b01100001;
DRAM[6534] = 8'b01101110;
DRAM[6535] = 8'b10001000;
DRAM[6536] = 8'b10011101;
DRAM[6537] = 8'b10101001;
DRAM[6538] = 8'b10101100;
DRAM[6539] = 8'b10101100;
DRAM[6540] = 8'b10101111;
DRAM[6541] = 8'b10101000;
DRAM[6542] = 8'b10010110;
DRAM[6543] = 8'b01110011;
DRAM[6544] = 8'b01001101;
DRAM[6545] = 8'b01001110;
DRAM[6546] = 8'b01010100;
DRAM[6547] = 8'b01011100;
DRAM[6548] = 8'b01011111;
DRAM[6549] = 8'b01100001;
DRAM[6550] = 8'b01100010;
DRAM[6551] = 8'b01100010;
DRAM[6552] = 8'b01100011;
DRAM[6553] = 8'b01011111;
DRAM[6554] = 8'b01100100;
DRAM[6555] = 8'b01101010;
DRAM[6556] = 8'b01101010;
DRAM[6557] = 8'b01101011;
DRAM[6558] = 8'b01100010;
DRAM[6559] = 8'b01011110;
DRAM[6560] = 8'b11010010;
DRAM[6561] = 8'b11000100;
DRAM[6562] = 8'b10111001;
DRAM[6563] = 8'b10100100;
DRAM[6564] = 8'b01111110;
DRAM[6565] = 8'b01111011;
DRAM[6566] = 8'b10000001;
DRAM[6567] = 8'b01110010;
DRAM[6568] = 8'b01111101;
DRAM[6569] = 8'b10000010;
DRAM[6570] = 8'b10000101;
DRAM[6571] = 8'b10000001;
DRAM[6572] = 8'b01111100;
DRAM[6573] = 8'b01111101;
DRAM[6574] = 8'b01111101;
DRAM[6575] = 8'b01100100;
DRAM[6576] = 8'b01011100;
DRAM[6577] = 8'b01001111;
DRAM[6578] = 8'b01001101;
DRAM[6579] = 8'b01010011;
DRAM[6580] = 8'b00110000;
DRAM[6581] = 8'b00100110;
DRAM[6582] = 8'b01001110;
DRAM[6583] = 8'b01010101;
DRAM[6584] = 8'b00101100;
DRAM[6585] = 8'b01000100;
DRAM[6586] = 8'b01010011;
DRAM[6587] = 8'b00110111;
DRAM[6588] = 8'b00110101;
DRAM[6589] = 8'b00110011;
DRAM[6590] = 8'b01010001;
DRAM[6591] = 8'b00110011;
DRAM[6592] = 8'b01110001;
DRAM[6593] = 8'b01110111;
DRAM[6594] = 8'b01110010;
DRAM[6595] = 8'b10010111;
DRAM[6596] = 8'b11000001;
DRAM[6597] = 8'b11000010;
DRAM[6598] = 8'b10111111;
DRAM[6599] = 8'b10110111;
DRAM[6600] = 8'b10110101;
DRAM[6601] = 8'b10110010;
DRAM[6602] = 8'b10110010;
DRAM[6603] = 8'b10101110;
DRAM[6604] = 8'b10101100;
DRAM[6605] = 8'b10110110;
DRAM[6606] = 8'b10110100;
DRAM[6607] = 8'b10111011;
DRAM[6608] = 8'b10110111;
DRAM[6609] = 8'b10111000;
DRAM[6610] = 8'b11000001;
DRAM[6611] = 8'b10101000;
DRAM[6612] = 8'b01100000;
DRAM[6613] = 8'b01010010;
DRAM[6614] = 8'b01101010;
DRAM[6615] = 8'b01100010;
DRAM[6616] = 8'b10000110;
DRAM[6617] = 8'b01110110;
DRAM[6618] = 8'b10010010;
DRAM[6619] = 8'b10101111;
DRAM[6620] = 8'b11000001;
DRAM[6621] = 8'b01110100;
DRAM[6622] = 8'b00101001;
DRAM[6623] = 8'b00101011;
DRAM[6624] = 8'b00101101;
DRAM[6625] = 8'b00110100;
DRAM[6626] = 8'b00110110;
DRAM[6627] = 8'b00110100;
DRAM[6628] = 8'b00110111;
DRAM[6629] = 8'b00110001;
DRAM[6630] = 8'b00101111;
DRAM[6631] = 8'b00110000;
DRAM[6632] = 8'b00111000;
DRAM[6633] = 8'b00111011;
DRAM[6634] = 8'b01100010;
DRAM[6635] = 8'b10000101;
DRAM[6636] = 8'b10000000;
DRAM[6637] = 8'b10011011;
DRAM[6638] = 8'b10101000;
DRAM[6639] = 8'b10100111;
DRAM[6640] = 8'b10100100;
DRAM[6641] = 8'b10100011;
DRAM[6642] = 8'b10100010;
DRAM[6643] = 8'b10100010;
DRAM[6644] = 8'b10100100;
DRAM[6645] = 8'b10100011;
DRAM[6646] = 8'b10100000;
DRAM[6647] = 8'b10011110;
DRAM[6648] = 8'b10100000;
DRAM[6649] = 8'b10011110;
DRAM[6650] = 8'b10011111;
DRAM[6651] = 8'b10011100;
DRAM[6652] = 8'b10011100;
DRAM[6653] = 8'b10011010;
DRAM[6654] = 8'b10011010;
DRAM[6655] = 8'b10010110;
DRAM[6656] = 8'b01101101;
DRAM[6657] = 8'b01101100;
DRAM[6658] = 8'b01101000;
DRAM[6659] = 8'b01100110;
DRAM[6660] = 8'b01100011;
DRAM[6661] = 8'b01100000;
DRAM[6662] = 8'b01101010;
DRAM[6663] = 8'b10001001;
DRAM[6664] = 8'b10011101;
DRAM[6665] = 8'b10101100;
DRAM[6666] = 8'b10101100;
DRAM[6667] = 8'b10101101;
DRAM[6668] = 8'b10101110;
DRAM[6669] = 8'b10100110;
DRAM[6670] = 8'b10010101;
DRAM[6671] = 8'b01110011;
DRAM[6672] = 8'b01001101;
DRAM[6673] = 8'b01001100;
DRAM[6674] = 8'b01010100;
DRAM[6675] = 8'b01011100;
DRAM[6676] = 8'b01011110;
DRAM[6677] = 8'b01100000;
DRAM[6678] = 8'b01100010;
DRAM[6679] = 8'b01011111;
DRAM[6680] = 8'b01100001;
DRAM[6681] = 8'b01100001;
DRAM[6682] = 8'b01100110;
DRAM[6683] = 8'b01101001;
DRAM[6684] = 8'b01101110;
DRAM[6685] = 8'b01101110;
DRAM[6686] = 8'b01101000;
DRAM[6687] = 8'b01011011;
DRAM[6688] = 8'b10011111;
DRAM[6689] = 8'b11001101;
DRAM[6690] = 8'b11000010;
DRAM[6691] = 8'b10100010;
DRAM[6692] = 8'b10001110;
DRAM[6693] = 8'b01110100;
DRAM[6694] = 8'b01110000;
DRAM[6695] = 8'b01111001;
DRAM[6696] = 8'b10000001;
DRAM[6697] = 8'b01110111;
DRAM[6698] = 8'b01110001;
DRAM[6699] = 8'b01111110;
DRAM[6700] = 8'b01111100;
DRAM[6701] = 8'b01111100;
DRAM[6702] = 8'b01100101;
DRAM[6703] = 8'b01001100;
DRAM[6704] = 8'b01000010;
DRAM[6705] = 8'b01010001;
DRAM[6706] = 8'b01011010;
DRAM[6707] = 8'b01001011;
DRAM[6708] = 8'b00110111;
DRAM[6709] = 8'b00101110;
DRAM[6710] = 8'b01010001;
DRAM[6711] = 8'b01001010;
DRAM[6712] = 8'b00111100;
DRAM[6713] = 8'b00111011;
DRAM[6714] = 8'b00110000;
DRAM[6715] = 8'b00111010;
DRAM[6716] = 8'b01001010;
DRAM[6717] = 8'b01001001;
DRAM[6718] = 8'b01010101;
DRAM[6719] = 8'b01001010;
DRAM[6720] = 8'b01100011;
DRAM[6721] = 8'b01111100;
DRAM[6722] = 8'b10001100;
DRAM[6723] = 8'b10101110;
DRAM[6724] = 8'b10110100;
DRAM[6725] = 8'b10110111;
DRAM[6726] = 8'b10111001;
DRAM[6727] = 8'b10110000;
DRAM[6728] = 8'b10101110;
DRAM[6729] = 8'b10101111;
DRAM[6730] = 8'b10101110;
DRAM[6731] = 8'b10101111;
DRAM[6732] = 8'b10101111;
DRAM[6733] = 8'b10110100;
DRAM[6734] = 8'b10110111;
DRAM[6735] = 8'b10111111;
DRAM[6736] = 8'b10111101;
DRAM[6737] = 8'b11000011;
DRAM[6738] = 8'b11001000;
DRAM[6739] = 8'b10111100;
DRAM[6740] = 8'b10000000;
DRAM[6741] = 8'b01010110;
DRAM[6742] = 8'b01001000;
DRAM[6743] = 8'b01011000;
DRAM[6744] = 8'b01011101;
DRAM[6745] = 8'b10000110;
DRAM[6746] = 8'b10001100;
DRAM[6747] = 8'b10011110;
DRAM[6748] = 8'b01011000;
DRAM[6749] = 8'b00101010;
DRAM[6750] = 8'b00101101;
DRAM[6751] = 8'b00101101;
DRAM[6752] = 8'b00101111;
DRAM[6753] = 8'b00110111;
DRAM[6754] = 8'b00111000;
DRAM[6755] = 8'b00111011;
DRAM[6756] = 8'b00110111;
DRAM[6757] = 8'b00101110;
DRAM[6758] = 8'b00110001;
DRAM[6759] = 8'b00110001;
DRAM[6760] = 8'b00110100;
DRAM[6761] = 8'b01000100;
DRAM[6762] = 8'b01111100;
DRAM[6763] = 8'b10000000;
DRAM[6764] = 8'b10000010;
DRAM[6765] = 8'b10100100;
DRAM[6766] = 8'b10101000;
DRAM[6767] = 8'b10101000;
DRAM[6768] = 8'b10100011;
DRAM[6769] = 8'b10100100;
DRAM[6770] = 8'b10100011;
DRAM[6771] = 8'b10100100;
DRAM[6772] = 8'b10100000;
DRAM[6773] = 8'b10100010;
DRAM[6774] = 8'b10100000;
DRAM[6775] = 8'b10100000;
DRAM[6776] = 8'b10100001;
DRAM[6777] = 8'b10011110;
DRAM[6778] = 8'b10011100;
DRAM[6779] = 8'b10011101;
DRAM[6780] = 8'b10011101;
DRAM[6781] = 8'b10011010;
DRAM[6782] = 8'b10011001;
DRAM[6783] = 8'b10010111;
DRAM[6784] = 8'b01101010;
DRAM[6785] = 8'b01101001;
DRAM[6786] = 8'b01101000;
DRAM[6787] = 8'b01100100;
DRAM[6788] = 8'b01100101;
DRAM[6789] = 8'b01011100;
DRAM[6790] = 8'b01101001;
DRAM[6791] = 8'b10000101;
DRAM[6792] = 8'b10011011;
DRAM[6793] = 8'b10101000;
DRAM[6794] = 8'b10101110;
DRAM[6795] = 8'b10101100;
DRAM[6796] = 8'b10101111;
DRAM[6797] = 8'b10101010;
DRAM[6798] = 8'b10010110;
DRAM[6799] = 8'b01110110;
DRAM[6800] = 8'b01001010;
DRAM[6801] = 8'b01001100;
DRAM[6802] = 8'b01010010;
DRAM[6803] = 8'b01011001;
DRAM[6804] = 8'b01011111;
DRAM[6805] = 8'b01100011;
DRAM[6806] = 8'b01100000;
DRAM[6807] = 8'b01100001;
DRAM[6808] = 8'b01100001;
DRAM[6809] = 8'b01100000;
DRAM[6810] = 8'b01100110;
DRAM[6811] = 8'b01101000;
DRAM[6812] = 8'b01101111;
DRAM[6813] = 8'b01101111;
DRAM[6814] = 8'b01101010;
DRAM[6815] = 8'b01011101;
DRAM[6816] = 8'b10011011;
DRAM[6817] = 8'b11010111;
DRAM[6818] = 8'b11001001;
DRAM[6819] = 8'b10101101;
DRAM[6820] = 8'b01111000;
DRAM[6821] = 8'b01111010;
DRAM[6822] = 8'b01101100;
DRAM[6823] = 8'b01111100;
DRAM[6824] = 8'b01110101;
DRAM[6825] = 8'b01111001;
DRAM[6826] = 8'b10001000;
DRAM[6827] = 8'b10000011;
DRAM[6828] = 8'b01101010;
DRAM[6829] = 8'b01111100;
DRAM[6830] = 8'b01011100;
DRAM[6831] = 8'b01000110;
DRAM[6832] = 8'b00111100;
DRAM[6833] = 8'b00110100;
DRAM[6834] = 8'b01001101;
DRAM[6835] = 8'b01000110;
DRAM[6836] = 8'b01000100;
DRAM[6837] = 8'b00111001;
DRAM[6838] = 8'b00111110;
DRAM[6839] = 8'b01101110;
DRAM[6840] = 8'b01000110;
DRAM[6841] = 8'b00101111;
DRAM[6842] = 8'b00101110;
DRAM[6843] = 8'b00110000;
DRAM[6844] = 8'b00110001;
DRAM[6845] = 8'b00101010;
DRAM[6846] = 8'b01000000;
DRAM[6847] = 8'b01100101;
DRAM[6848] = 8'b01001011;
DRAM[6849] = 8'b10000101;
DRAM[6850] = 8'b10100001;
DRAM[6851] = 8'b10101110;
DRAM[6852] = 8'b10110010;
DRAM[6853] = 8'b10110110;
DRAM[6854] = 8'b10101101;
DRAM[6855] = 8'b10101001;
DRAM[6856] = 8'b10110000;
DRAM[6857] = 8'b10101110;
DRAM[6858] = 8'b10101111;
DRAM[6859] = 8'b10101101;
DRAM[6860] = 8'b10101011;
DRAM[6861] = 8'b10111000;
DRAM[6862] = 8'b11000110;
DRAM[6863] = 8'b11000101;
DRAM[6864] = 8'b11000100;
DRAM[6865] = 8'b11000100;
DRAM[6866] = 8'b11000110;
DRAM[6867] = 8'b11000011;
DRAM[6868] = 8'b10011101;
DRAM[6869] = 8'b01100100;
DRAM[6870] = 8'b01000010;
DRAM[6871] = 8'b01000100;
DRAM[6872] = 8'b01001110;
DRAM[6873] = 8'b01111101;
DRAM[6874] = 8'b10010000;
DRAM[6875] = 8'b10001010;
DRAM[6876] = 8'b01001100;
DRAM[6877] = 8'b00101011;
DRAM[6878] = 8'b00101001;
DRAM[6879] = 8'b00101011;
DRAM[6880] = 8'b00111000;
DRAM[6881] = 8'b00110101;
DRAM[6882] = 8'b00111011;
DRAM[6883] = 8'b00111010;
DRAM[6884] = 8'b00110000;
DRAM[6885] = 8'b00101011;
DRAM[6886] = 8'b00101101;
DRAM[6887] = 8'b00110101;
DRAM[6888] = 8'b00110110;
DRAM[6889] = 8'b01010111;
DRAM[6890] = 8'b10000110;
DRAM[6891] = 8'b01111101;
DRAM[6892] = 8'b10001110;
DRAM[6893] = 8'b10100010;
DRAM[6894] = 8'b10100101;
DRAM[6895] = 8'b10100110;
DRAM[6896] = 8'b10100111;
DRAM[6897] = 8'b10100100;
DRAM[6898] = 8'b10100010;
DRAM[6899] = 8'b10100100;
DRAM[6900] = 8'b10100000;
DRAM[6901] = 8'b10100011;
DRAM[6902] = 8'b10100010;
DRAM[6903] = 8'b10100010;
DRAM[6904] = 8'b10100010;
DRAM[6905] = 8'b10011111;
DRAM[6906] = 8'b10011110;
DRAM[6907] = 8'b10011101;
DRAM[6908] = 8'b10011100;
DRAM[6909] = 8'b10011100;
DRAM[6910] = 8'b10011010;
DRAM[6911] = 8'b10011000;
DRAM[6912] = 8'b01101010;
DRAM[6913] = 8'b01101001;
DRAM[6914] = 8'b01101001;
DRAM[6915] = 8'b01100100;
DRAM[6916] = 8'b01100001;
DRAM[6917] = 8'b01011001;
DRAM[6918] = 8'b01100100;
DRAM[6919] = 8'b10001000;
DRAM[6920] = 8'b10011001;
DRAM[6921] = 8'b10101001;
DRAM[6922] = 8'b10101100;
DRAM[6923] = 8'b10101101;
DRAM[6924] = 8'b10101110;
DRAM[6925] = 8'b10100111;
DRAM[6926] = 8'b10010110;
DRAM[6927] = 8'b01110110;
DRAM[6928] = 8'b01001100;
DRAM[6929] = 8'b01001010;
DRAM[6930] = 8'b01011001;
DRAM[6931] = 8'b01011101;
DRAM[6932] = 8'b01100001;
DRAM[6933] = 8'b01100010;
DRAM[6934] = 8'b01100110;
DRAM[6935] = 8'b01100110;
DRAM[6936] = 8'b01100011;
DRAM[6937] = 8'b01100010;
DRAM[6938] = 8'b01100101;
DRAM[6939] = 8'b01101011;
DRAM[6940] = 8'b01110000;
DRAM[6941] = 8'b01110000;
DRAM[6942] = 8'b01101100;
DRAM[6943] = 8'b01100100;
DRAM[6944] = 8'b10010110;
DRAM[6945] = 8'b11010110;
DRAM[6946] = 8'b11010100;
DRAM[6947] = 8'b01111001;
DRAM[6948] = 8'b01110010;
DRAM[6949] = 8'b01110100;
DRAM[6950] = 8'b01111001;
DRAM[6951] = 8'b01110011;
DRAM[6952] = 8'b01110110;
DRAM[6953] = 8'b10000111;
DRAM[6954] = 8'b10000100;
DRAM[6955] = 8'b01111100;
DRAM[6956] = 8'b01011001;
DRAM[6957] = 8'b00111100;
DRAM[6958] = 8'b00111110;
DRAM[6959] = 8'b01000010;
DRAM[6960] = 8'b00101101;
DRAM[6961] = 8'b00110000;
DRAM[6962] = 8'b01000110;
DRAM[6963] = 8'b01000100;
DRAM[6964] = 8'b01011001;
DRAM[6965] = 8'b00101100;
DRAM[6966] = 8'b00111010;
DRAM[6967] = 8'b01001111;
DRAM[6968] = 8'b01110111;
DRAM[6969] = 8'b00110011;
DRAM[6970] = 8'b00101111;
DRAM[6971] = 8'b00101000;
DRAM[6972] = 8'b00100111;
DRAM[6973] = 8'b00110100;
DRAM[6974] = 8'b01110100;
DRAM[6975] = 8'b01100100;
DRAM[6976] = 8'b10001011;
DRAM[6977] = 8'b10100011;
DRAM[6978] = 8'b10110101;
DRAM[6979] = 8'b10110111;
DRAM[6980] = 8'b10111101;
DRAM[6981] = 8'b10110101;
DRAM[6982] = 8'b10100010;
DRAM[6983] = 8'b10100100;
DRAM[6984] = 8'b10101011;
DRAM[6985] = 8'b10110011;
DRAM[6986] = 8'b10100001;
DRAM[6987] = 8'b10101100;
DRAM[6988] = 8'b10110111;
DRAM[6989] = 8'b11000010;
DRAM[6990] = 8'b11000101;
DRAM[6991] = 8'b11001000;
DRAM[6992] = 8'b11000100;
DRAM[6993] = 8'b11000111;
DRAM[6994] = 8'b11001010;
DRAM[6995] = 8'b11000100;
DRAM[6996] = 8'b10101010;
DRAM[6997] = 8'b01101010;
DRAM[6998] = 8'b01000010;
DRAM[6999] = 8'b00101110;
DRAM[7000] = 8'b01010010;
DRAM[7001] = 8'b01100110;
DRAM[7002] = 8'b10001111;
DRAM[7003] = 8'b10010011;
DRAM[7004] = 8'b00111100;
DRAM[7005] = 8'b00101110;
DRAM[7006] = 8'b00101101;
DRAM[7007] = 8'b00101111;
DRAM[7008] = 8'b00110111;
DRAM[7009] = 8'b00110111;
DRAM[7010] = 8'b00111101;
DRAM[7011] = 8'b00111010;
DRAM[7012] = 8'b00110010;
DRAM[7013] = 8'b00101010;
DRAM[7014] = 8'b00110100;
DRAM[7015] = 8'b00101101;
DRAM[7016] = 8'b00110111;
DRAM[7017] = 8'b01110110;
DRAM[7018] = 8'b10001000;
DRAM[7019] = 8'b10000010;
DRAM[7020] = 8'b10010111;
DRAM[7021] = 8'b10011101;
DRAM[7022] = 8'b10100100;
DRAM[7023] = 8'b10100101;
DRAM[7024] = 8'b10100100;
DRAM[7025] = 8'b10100011;
DRAM[7026] = 8'b10100001;
DRAM[7027] = 8'b10100000;
DRAM[7028] = 8'b10100001;
DRAM[7029] = 8'b10100100;
DRAM[7030] = 8'b10100010;
DRAM[7031] = 8'b10100000;
DRAM[7032] = 8'b10011111;
DRAM[7033] = 8'b10011111;
DRAM[7034] = 8'b10011101;
DRAM[7035] = 8'b10011110;
DRAM[7036] = 8'b10011110;
DRAM[7037] = 8'b10011011;
DRAM[7038] = 8'b10011010;
DRAM[7039] = 8'b10010101;
DRAM[7040] = 8'b01100111;
DRAM[7041] = 8'b01101100;
DRAM[7042] = 8'b01100110;
DRAM[7043] = 8'b01100011;
DRAM[7044] = 8'b01100100;
DRAM[7045] = 8'b01011100;
DRAM[7046] = 8'b01101000;
DRAM[7047] = 8'b10000111;
DRAM[7048] = 8'b10011011;
DRAM[7049] = 8'b10101001;
DRAM[7050] = 8'b10101100;
DRAM[7051] = 8'b10101110;
DRAM[7052] = 8'b10101101;
DRAM[7053] = 8'b10101000;
DRAM[7054] = 8'b10011000;
DRAM[7055] = 8'b01110101;
DRAM[7056] = 8'b01010000;
DRAM[7057] = 8'b01001010;
DRAM[7058] = 8'b01010100;
DRAM[7059] = 8'b01100000;
DRAM[7060] = 8'b01100100;
DRAM[7061] = 8'b01100001;
DRAM[7062] = 8'b01100100;
DRAM[7063] = 8'b01100011;
DRAM[7064] = 8'b01100100;
DRAM[7065] = 8'b01100101;
DRAM[7066] = 8'b01100110;
DRAM[7067] = 8'b01101010;
DRAM[7068] = 8'b01101101;
DRAM[7069] = 8'b01110100;
DRAM[7070] = 8'b01101111;
DRAM[7071] = 8'b01101010;
DRAM[7072] = 8'b01110101;
DRAM[7073] = 8'b11011011;
DRAM[7074] = 8'b10111000;
DRAM[7075] = 8'b01101010;
DRAM[7076] = 8'b01101010;
DRAM[7077] = 8'b01110010;
DRAM[7078] = 8'b01101111;
DRAM[7079] = 8'b01111010;
DRAM[7080] = 8'b01111111;
DRAM[7081] = 8'b01101110;
DRAM[7082] = 8'b01110110;
DRAM[7083] = 8'b01101110;
DRAM[7084] = 8'b01011001;
DRAM[7085] = 8'b00101110;
DRAM[7086] = 8'b01010011;
DRAM[7087] = 8'b00101010;
DRAM[7088] = 8'b00110000;
DRAM[7089] = 8'b00110001;
DRAM[7090] = 8'b00110011;
DRAM[7091] = 8'b01001011;
DRAM[7092] = 8'b01000111;
DRAM[7093] = 8'b00111010;
DRAM[7094] = 8'b01000011;
DRAM[7095] = 8'b00110010;
DRAM[7096] = 8'b01110101;
DRAM[7097] = 8'b01000010;
DRAM[7098] = 8'b00111001;
DRAM[7099] = 8'b00100010;
DRAM[7100] = 8'b00101010;
DRAM[7101] = 8'b10001000;
DRAM[7102] = 8'b01110011;
DRAM[7103] = 8'b10100101;
DRAM[7104] = 8'b10011110;
DRAM[7105] = 8'b10010011;
DRAM[7106] = 8'b10110010;
DRAM[7107] = 8'b10111010;
DRAM[7108] = 8'b10111100;
DRAM[7109] = 8'b10101001;
DRAM[7110] = 8'b10100100;
DRAM[7111] = 8'b10100110;
DRAM[7112] = 8'b10110100;
DRAM[7113] = 8'b10100010;
DRAM[7114] = 8'b10100110;
DRAM[7115] = 8'b10110001;
DRAM[7116] = 8'b10111100;
DRAM[7117] = 8'b11000100;
DRAM[7118] = 8'b11000110;
DRAM[7119] = 8'b11001100;
DRAM[7120] = 8'b11001010;
DRAM[7121] = 8'b11001101;
DRAM[7122] = 8'b11010000;
DRAM[7123] = 8'b11001110;
DRAM[7124] = 8'b10111000;
DRAM[7125] = 8'b01111100;
DRAM[7126] = 8'b01001011;
DRAM[7127] = 8'b00101001;
DRAM[7128] = 8'b00111101;
DRAM[7129] = 8'b01010100;
DRAM[7130] = 8'b10011100;
DRAM[7131] = 8'b10001110;
DRAM[7132] = 8'b00110001;
DRAM[7133] = 8'b00101100;
DRAM[7134] = 8'b00110000;
DRAM[7135] = 8'b00110011;
DRAM[7136] = 8'b00110110;
DRAM[7137] = 8'b00110110;
DRAM[7138] = 8'b00111110;
DRAM[7139] = 8'b00110110;
DRAM[7140] = 8'b00101011;
DRAM[7141] = 8'b00101100;
DRAM[7142] = 8'b00110011;
DRAM[7143] = 8'b00110101;
DRAM[7144] = 8'b01010001;
DRAM[7145] = 8'b10001010;
DRAM[7146] = 8'b10000100;
DRAM[7147] = 8'b10010000;
DRAM[7148] = 8'b10011000;
DRAM[7149] = 8'b10010110;
DRAM[7150] = 8'b10011011;
DRAM[7151] = 8'b10011101;
DRAM[7152] = 8'b10100001;
DRAM[7153] = 8'b10100011;
DRAM[7154] = 8'b10100000;
DRAM[7155] = 8'b10100001;
DRAM[7156] = 8'b10100000;
DRAM[7157] = 8'b10100000;
DRAM[7158] = 8'b10100101;
DRAM[7159] = 8'b10100000;
DRAM[7160] = 8'b10100000;
DRAM[7161] = 8'b10011101;
DRAM[7162] = 8'b10011110;
DRAM[7163] = 8'b10011110;
DRAM[7164] = 8'b10011110;
DRAM[7165] = 8'b10011011;
DRAM[7166] = 8'b10011010;
DRAM[7167] = 8'b10011000;
DRAM[7168] = 8'b01100111;
DRAM[7169] = 8'b01100110;
DRAM[7170] = 8'b01100110;
DRAM[7171] = 8'b01100011;
DRAM[7172] = 8'b01100010;
DRAM[7173] = 8'b01011100;
DRAM[7174] = 8'b01100011;
DRAM[7175] = 8'b10000111;
DRAM[7176] = 8'b10011011;
DRAM[7177] = 8'b10100111;
DRAM[7178] = 8'b10101100;
DRAM[7179] = 8'b10101110;
DRAM[7180] = 8'b10101101;
DRAM[7181] = 8'b10101011;
DRAM[7182] = 8'b10010110;
DRAM[7183] = 8'b01111010;
DRAM[7184] = 8'b01010001;
DRAM[7185] = 8'b01001110;
DRAM[7186] = 8'b01010100;
DRAM[7187] = 8'b01011110;
DRAM[7188] = 8'b01100100;
DRAM[7189] = 8'b01100101;
DRAM[7190] = 8'b01101000;
DRAM[7191] = 8'b01100110;
DRAM[7192] = 8'b01100100;
DRAM[7193] = 8'b01100011;
DRAM[7194] = 8'b01100110;
DRAM[7195] = 8'b01111001;
DRAM[7196] = 8'b01111111;
DRAM[7197] = 8'b01110011;
DRAM[7198] = 8'b01110010;
DRAM[7199] = 8'b01101110;
DRAM[7200] = 8'b01100100;
DRAM[7201] = 8'b11001110;
DRAM[7202] = 8'b10100010;
DRAM[7203] = 8'b01110011;
DRAM[7204] = 8'b01111000;
DRAM[7205] = 8'b01101011;
DRAM[7206] = 8'b01110110;
DRAM[7207] = 8'b01111110;
DRAM[7208] = 8'b01111000;
DRAM[7209] = 8'b01100100;
DRAM[7210] = 8'b01001000;
DRAM[7211] = 8'b01000100;
DRAM[7212] = 8'b01001001;
DRAM[7213] = 8'b00110101;
DRAM[7214] = 8'b01001100;
DRAM[7215] = 8'b00101010;
DRAM[7216] = 8'b00111011;
DRAM[7217] = 8'b00110100;
DRAM[7218] = 8'b00110010;
DRAM[7219] = 8'b00110110;
DRAM[7220] = 8'b01000000;
DRAM[7221] = 8'b00111001;
DRAM[7222] = 8'b01010111;
DRAM[7223] = 8'b01010011;
DRAM[7224] = 8'b01100010;
DRAM[7225] = 8'b00101001;
DRAM[7226] = 8'b00100010;
DRAM[7227] = 8'b00011101;
DRAM[7228] = 8'b01111101;
DRAM[7229] = 8'b01110110;
DRAM[7230] = 8'b10100100;
DRAM[7231] = 8'b10101011;
DRAM[7232] = 8'b10100101;
DRAM[7233] = 8'b10010111;
DRAM[7234] = 8'b10100111;
DRAM[7235] = 8'b10111010;
DRAM[7236] = 8'b10110010;
DRAM[7237] = 8'b10101010;
DRAM[7238] = 8'b10101011;
DRAM[7239] = 8'b10101010;
DRAM[7240] = 8'b10011010;
DRAM[7241] = 8'b10100100;
DRAM[7242] = 8'b10101101;
DRAM[7243] = 8'b10111001;
DRAM[7244] = 8'b10111110;
DRAM[7245] = 8'b11000100;
DRAM[7246] = 8'b11000110;
DRAM[7247] = 8'b11001001;
DRAM[7248] = 8'b11001001;
DRAM[7249] = 8'b11001110;
DRAM[7250] = 8'b11010001;
DRAM[7251] = 8'b11010010;
DRAM[7252] = 8'b11000100;
DRAM[7253] = 8'b10001101;
DRAM[7254] = 8'b01010101;
DRAM[7255] = 8'b00101111;
DRAM[7256] = 8'b00101011;
DRAM[7257] = 8'b01000000;
DRAM[7258] = 8'b10010101;
DRAM[7259] = 8'b10011100;
DRAM[7260] = 8'b00110100;
DRAM[7261] = 8'b00110101;
DRAM[7262] = 8'b00110001;
DRAM[7263] = 8'b00111000;
DRAM[7264] = 8'b00110110;
DRAM[7265] = 8'b00111110;
DRAM[7266] = 8'b01000000;
DRAM[7267] = 8'b00110001;
DRAM[7268] = 8'b00101110;
DRAM[7269] = 8'b00110011;
DRAM[7270] = 8'b00110101;
DRAM[7271] = 8'b00101100;
DRAM[7272] = 8'b01101011;
DRAM[7273] = 8'b10001101;
DRAM[7274] = 8'b10000011;
DRAM[7275] = 8'b10011101;
DRAM[7276] = 8'b10011100;
DRAM[7277] = 8'b10010111;
DRAM[7278] = 8'b10010110;
DRAM[7279] = 8'b10010110;
DRAM[7280] = 8'b10010111;
DRAM[7281] = 8'b10010111;
DRAM[7282] = 8'b10011100;
DRAM[7283] = 8'b10011110;
DRAM[7284] = 8'b10011111;
DRAM[7285] = 8'b10011111;
DRAM[7286] = 8'b10100001;
DRAM[7287] = 8'b10100001;
DRAM[7288] = 8'b10011111;
DRAM[7289] = 8'b10100000;
DRAM[7290] = 8'b10011111;
DRAM[7291] = 8'b10011100;
DRAM[7292] = 8'b10011100;
DRAM[7293] = 8'b10011010;
DRAM[7294] = 8'b10011100;
DRAM[7295] = 8'b10010111;
DRAM[7296] = 8'b01101001;
DRAM[7297] = 8'b01101000;
DRAM[7298] = 8'b01100100;
DRAM[7299] = 8'b01100100;
DRAM[7300] = 8'b01100010;
DRAM[7301] = 8'b01011100;
DRAM[7302] = 8'b01100111;
DRAM[7303] = 8'b10000101;
DRAM[7304] = 8'b10011001;
DRAM[7305] = 8'b10101011;
DRAM[7306] = 8'b10101100;
DRAM[7307] = 8'b10101110;
DRAM[7308] = 8'b10101101;
DRAM[7309] = 8'b10101001;
DRAM[7310] = 8'b10010100;
DRAM[7311] = 8'b01111000;
DRAM[7312] = 8'b01010011;
DRAM[7313] = 8'b01010000;
DRAM[7314] = 8'b01010111;
DRAM[7315] = 8'b01100011;
DRAM[7316] = 8'b01100110;
DRAM[7317] = 8'b01100101;
DRAM[7318] = 8'b01101000;
DRAM[7319] = 8'b01100110;
DRAM[7320] = 8'b01100100;
DRAM[7321] = 8'b01100101;
DRAM[7322] = 8'b01101000;
DRAM[7323] = 8'b01111000;
DRAM[7324] = 8'b01110011;
DRAM[7325] = 8'b01110100;
DRAM[7326] = 8'b01110110;
DRAM[7327] = 8'b01110100;
DRAM[7328] = 8'b01101111;
DRAM[7329] = 8'b10011000;
DRAM[7330] = 8'b10110010;
DRAM[7331] = 8'b01110101;
DRAM[7332] = 8'b01110000;
DRAM[7333] = 8'b01111100;
DRAM[7334] = 8'b01111100;
DRAM[7335] = 8'b10000001;
DRAM[7336] = 8'b01111100;
DRAM[7337] = 8'b01100101;
DRAM[7338] = 8'b01000110;
DRAM[7339] = 8'b00111011;
DRAM[7340] = 8'b00101100;
DRAM[7341] = 8'b00101101;
DRAM[7342] = 8'b01001010;
DRAM[7343] = 8'b00110010;
DRAM[7344] = 8'b00111001;
DRAM[7345] = 8'b00110111;
DRAM[7346] = 8'b00110100;
DRAM[7347] = 8'b00110010;
DRAM[7348] = 8'b00111100;
DRAM[7349] = 8'b00110101;
DRAM[7350] = 8'b01011100;
DRAM[7351] = 8'b01011100;
DRAM[7352] = 8'b01011010;
DRAM[7353] = 8'b01001010;
DRAM[7354] = 8'b00011110;
DRAM[7355] = 8'b01110000;
DRAM[7356] = 8'b10000001;
DRAM[7357] = 8'b10100110;
DRAM[7358] = 8'b10101111;
DRAM[7359] = 8'b10110100;
DRAM[7360] = 8'b10101110;
DRAM[7361] = 8'b10010110;
DRAM[7362] = 8'b10101010;
DRAM[7363] = 8'b11000010;
DRAM[7364] = 8'b10110001;
DRAM[7365] = 8'b10100111;
DRAM[7366] = 8'b10100000;
DRAM[7367] = 8'b10011000;
DRAM[7368] = 8'b10011111;
DRAM[7369] = 8'b10101001;
DRAM[7370] = 8'b10110001;
DRAM[7371] = 8'b10111100;
DRAM[7372] = 8'b11000010;
DRAM[7373] = 8'b11000100;
DRAM[7374] = 8'b11000111;
DRAM[7375] = 8'b11001011;
DRAM[7376] = 8'b11001011;
DRAM[7377] = 8'b11010001;
DRAM[7378] = 8'b11010010;
DRAM[7379] = 8'b11010100;
DRAM[7380] = 8'b11001010;
DRAM[7381] = 8'b10011101;
DRAM[7382] = 8'b01011101;
DRAM[7383] = 8'b00110010;
DRAM[7384] = 8'b00100101;
DRAM[7385] = 8'b01000010;
DRAM[7386] = 8'b01101110;
DRAM[7387] = 8'b10010010;
DRAM[7388] = 8'b01000100;
DRAM[7389] = 8'b00110101;
DRAM[7390] = 8'b00110110;
DRAM[7391] = 8'b00110111;
DRAM[7392] = 8'b00111110;
DRAM[7393] = 8'b00111100;
DRAM[7394] = 8'b00111111;
DRAM[7395] = 8'b00110000;
DRAM[7396] = 8'b00101100;
DRAM[7397] = 8'b00110010;
DRAM[7398] = 8'b00101110;
DRAM[7399] = 8'b00111001;
DRAM[7400] = 8'b10000001;
DRAM[7401] = 8'b10001010;
DRAM[7402] = 8'b10001101;
DRAM[7403] = 8'b10100011;
DRAM[7404] = 8'b10100001;
DRAM[7405] = 8'b10011101;
DRAM[7406] = 8'b10011011;
DRAM[7407] = 8'b10011000;
DRAM[7408] = 8'b10010101;
DRAM[7409] = 8'b10010100;
DRAM[7410] = 8'b10011000;
DRAM[7411] = 8'b10010101;
DRAM[7412] = 8'b10010101;
DRAM[7413] = 8'b10011001;
DRAM[7414] = 8'b10011101;
DRAM[7415] = 8'b10011110;
DRAM[7416] = 8'b10011110;
DRAM[7417] = 8'b10011101;
DRAM[7418] = 8'b10011100;
DRAM[7419] = 8'b10011011;
DRAM[7420] = 8'b10011011;
DRAM[7421] = 8'b10011001;
DRAM[7422] = 8'b10011000;
DRAM[7423] = 8'b10010101;
DRAM[7424] = 8'b01100111;
DRAM[7425] = 8'b01100101;
DRAM[7426] = 8'b01100110;
DRAM[7427] = 8'b01100001;
DRAM[7428] = 8'b01011110;
DRAM[7429] = 8'b01011010;
DRAM[7430] = 8'b01100101;
DRAM[7431] = 8'b10000101;
DRAM[7432] = 8'b10011010;
DRAM[7433] = 8'b10101000;
DRAM[7434] = 8'b10101101;
DRAM[7435] = 8'b10110001;
DRAM[7436] = 8'b10101100;
DRAM[7437] = 8'b10101010;
DRAM[7438] = 8'b10010111;
DRAM[7439] = 8'b01110111;
DRAM[7440] = 8'b01010000;
DRAM[7441] = 8'b01010000;
DRAM[7442] = 8'b01011101;
DRAM[7443] = 8'b01011110;
DRAM[7444] = 8'b01100010;
DRAM[7445] = 8'b01100111;
DRAM[7446] = 8'b01101001;
DRAM[7447] = 8'b01100110;
DRAM[7448] = 8'b01100100;
DRAM[7449] = 8'b01101000;
DRAM[7450] = 8'b01101001;
DRAM[7451] = 8'b01110110;
DRAM[7452] = 8'b01110010;
DRAM[7453] = 8'b01111000;
DRAM[7454] = 8'b01110111;
DRAM[7455] = 8'b01111000;
DRAM[7456] = 8'b01110100;
DRAM[7457] = 8'b01110101;
DRAM[7458] = 8'b10110001;
DRAM[7459] = 8'b01111000;
DRAM[7460] = 8'b01111000;
DRAM[7461] = 8'b10000001;
DRAM[7462] = 8'b10000010;
DRAM[7463] = 8'b10000010;
DRAM[7464] = 8'b01011100;
DRAM[7465] = 8'b00111101;
DRAM[7466] = 8'b00110100;
DRAM[7467] = 8'b01010000;
DRAM[7468] = 8'b00101101;
DRAM[7469] = 8'b00101001;
DRAM[7470] = 8'b01010000;
DRAM[7471] = 8'b00110111;
DRAM[7472] = 8'b01000100;
DRAM[7473] = 8'b00110011;
DRAM[7474] = 8'b00110000;
DRAM[7475] = 8'b00111011;
DRAM[7476] = 8'b00111110;
DRAM[7477] = 8'b00101110;
DRAM[7478] = 8'b01001011;
DRAM[7479] = 8'b00111010;
DRAM[7480] = 8'b00011110;
DRAM[7481] = 8'b01100010;
DRAM[7482] = 8'b01100010;
DRAM[7483] = 8'b10000010;
DRAM[7484] = 8'b10001101;
DRAM[7485] = 8'b10100110;
DRAM[7486] = 8'b10110001;
DRAM[7487] = 8'b10111100;
DRAM[7488] = 8'b10110100;
DRAM[7489] = 8'b10001110;
DRAM[7490] = 8'b10110000;
DRAM[7491] = 8'b10111011;
DRAM[7492] = 8'b10100010;
DRAM[7493] = 8'b10100001;
DRAM[7494] = 8'b10011101;
DRAM[7495] = 8'b10011110;
DRAM[7496] = 8'b10101010;
DRAM[7497] = 8'b10101111;
DRAM[7498] = 8'b10110001;
DRAM[7499] = 8'b10111010;
DRAM[7500] = 8'b11000011;
DRAM[7501] = 8'b11000100;
DRAM[7502] = 8'b11000111;
DRAM[7503] = 8'b11001010;
DRAM[7504] = 8'b11001101;
DRAM[7505] = 8'b11010000;
DRAM[7506] = 8'b11010010;
DRAM[7507] = 8'b11010100;
DRAM[7508] = 8'b11010001;
DRAM[7509] = 8'b10101101;
DRAM[7510] = 8'b01101101;
DRAM[7511] = 8'b00111111;
DRAM[7512] = 8'b00101010;
DRAM[7513] = 8'b00101110;
DRAM[7514] = 8'b01110101;
DRAM[7515] = 8'b10100100;
DRAM[7516] = 8'b01010010;
DRAM[7517] = 8'b00110000;
DRAM[7518] = 8'b00110111;
DRAM[7519] = 8'b00111001;
DRAM[7520] = 8'b00111100;
DRAM[7521] = 8'b00111011;
DRAM[7522] = 8'b00111100;
DRAM[7523] = 8'b00110100;
DRAM[7524] = 8'b00110010;
DRAM[7525] = 8'b00110101;
DRAM[7526] = 8'b00101011;
DRAM[7527] = 8'b01010101;
DRAM[7528] = 8'b10001110;
DRAM[7529] = 8'b10000101;
DRAM[7530] = 8'b10010111;
DRAM[7531] = 8'b10100110;
DRAM[7532] = 8'b10100010;
DRAM[7533] = 8'b10100011;
DRAM[7534] = 8'b10100001;
DRAM[7535] = 8'b10100000;
DRAM[7536] = 8'b10011010;
DRAM[7537] = 8'b10011001;
DRAM[7538] = 8'b10011000;
DRAM[7539] = 8'b10010111;
DRAM[7540] = 8'b10010001;
DRAM[7541] = 8'b10010001;
DRAM[7542] = 8'b10010010;
DRAM[7543] = 8'b10010100;
DRAM[7544] = 8'b10010101;
DRAM[7545] = 8'b10010111;
DRAM[7546] = 8'b10011010;
DRAM[7547] = 8'b10011001;
DRAM[7548] = 8'b10010111;
DRAM[7549] = 8'b10011011;
DRAM[7550] = 8'b10011001;
DRAM[7551] = 8'b10011000;
DRAM[7552] = 8'b01101000;
DRAM[7553] = 8'b01100110;
DRAM[7554] = 8'b01100110;
DRAM[7555] = 8'b01100000;
DRAM[7556] = 8'b01100100;
DRAM[7557] = 8'b01011100;
DRAM[7558] = 8'b01100110;
DRAM[7559] = 8'b10000011;
DRAM[7560] = 8'b10011000;
DRAM[7561] = 8'b10101001;
DRAM[7562] = 8'b10101110;
DRAM[7563] = 8'b10101110;
DRAM[7564] = 8'b10101111;
DRAM[7565] = 8'b10101000;
DRAM[7566] = 8'b10011000;
DRAM[7567] = 8'b01110110;
DRAM[7568] = 8'b01010001;
DRAM[7569] = 8'b01001110;
DRAM[7570] = 8'b01010111;
DRAM[7571] = 8'b01011111;
DRAM[7572] = 8'b01100011;
DRAM[7573] = 8'b01100110;
DRAM[7574] = 8'b01100111;
DRAM[7575] = 8'b01100111;
DRAM[7576] = 8'b01100101;
DRAM[7577] = 8'b01100110;
DRAM[7578] = 8'b01101011;
DRAM[7579] = 8'b01110001;
DRAM[7580] = 8'b01110101;
DRAM[7581] = 8'b01110100;
DRAM[7582] = 8'b01110011;
DRAM[7583] = 8'b01101111;
DRAM[7584] = 8'b01110100;
DRAM[7585] = 8'b01111010;
DRAM[7586] = 8'b01101111;
DRAM[7587] = 8'b01110001;
DRAM[7588] = 8'b10000001;
DRAM[7589] = 8'b10000111;
DRAM[7590] = 8'b01111110;
DRAM[7591] = 8'b01101110;
DRAM[7592] = 8'b00111100;
DRAM[7593] = 8'b01000000;
DRAM[7594] = 8'b00100010;
DRAM[7595] = 8'b01011011;
DRAM[7596] = 8'b00111000;
DRAM[7597] = 8'b00110010;
DRAM[7598] = 8'b00101110;
DRAM[7599] = 8'b01000100;
DRAM[7600] = 8'b01000110;
DRAM[7601] = 8'b00100111;
DRAM[7602] = 8'b00101111;
DRAM[7603] = 8'b01001110;
DRAM[7604] = 8'b00111011;
DRAM[7605] = 8'b00111101;
DRAM[7606] = 8'b00110000;
DRAM[7607] = 8'b01010010;
DRAM[7608] = 8'b00011111;
DRAM[7609] = 8'b01001001;
DRAM[7610] = 8'b01111101;
DRAM[7611] = 8'b10001001;
DRAM[7612] = 8'b10100101;
DRAM[7613] = 8'b10100001;
DRAM[7614] = 8'b10101010;
DRAM[7615] = 8'b10111011;
DRAM[7616] = 8'b10111000;
DRAM[7617] = 8'b10011100;
DRAM[7618] = 8'b10110101;
DRAM[7619] = 8'b10101000;
DRAM[7620] = 8'b10011011;
DRAM[7621] = 8'b10100000;
DRAM[7622] = 8'b10100001;
DRAM[7623] = 8'b10100101;
DRAM[7624] = 8'b10101100;
DRAM[7625] = 8'b10101110;
DRAM[7626] = 8'b10110010;
DRAM[7627] = 8'b10110111;
DRAM[7628] = 8'b11000000;
DRAM[7629] = 8'b11000101;
DRAM[7630] = 8'b11000111;
DRAM[7631] = 8'b11000111;
DRAM[7632] = 8'b11001010;
DRAM[7633] = 8'b11001110;
DRAM[7634] = 8'b11010000;
DRAM[7635] = 8'b11010100;
DRAM[7636] = 8'b11010010;
DRAM[7637] = 8'b10111100;
DRAM[7638] = 8'b01110110;
DRAM[7639] = 8'b01001110;
DRAM[7640] = 8'b00101001;
DRAM[7641] = 8'b00101100;
DRAM[7642] = 8'b01011101;
DRAM[7643] = 8'b10110000;
DRAM[7644] = 8'b01000100;
DRAM[7645] = 8'b00110011;
DRAM[7646] = 8'b00111001;
DRAM[7647] = 8'b00111011;
DRAM[7648] = 8'b00111101;
DRAM[7649] = 8'b01000000;
DRAM[7650] = 8'b00110100;
DRAM[7651] = 8'b00110010;
DRAM[7652] = 8'b00110101;
DRAM[7653] = 8'b00110011;
DRAM[7654] = 8'b00111010;
DRAM[7655] = 8'b01111101;
DRAM[7656] = 8'b10001011;
DRAM[7657] = 8'b10001011;
DRAM[7658] = 8'b10100000;
DRAM[7659] = 8'b10100011;
DRAM[7660] = 8'b10100001;
DRAM[7661] = 8'b10100001;
DRAM[7662] = 8'b10100000;
DRAM[7663] = 8'b10100011;
DRAM[7664] = 8'b10100011;
DRAM[7665] = 8'b10100010;
DRAM[7666] = 8'b10011101;
DRAM[7667] = 8'b10011100;
DRAM[7668] = 8'b10010101;
DRAM[7669] = 8'b10010011;
DRAM[7670] = 8'b10010010;
DRAM[7671] = 8'b10010001;
DRAM[7672] = 8'b10001111;
DRAM[7673] = 8'b10001110;
DRAM[7674] = 8'b10010001;
DRAM[7675] = 8'b10010010;
DRAM[7676] = 8'b10010110;
DRAM[7677] = 8'b10011001;
DRAM[7678] = 8'b10010111;
DRAM[7679] = 8'b10010111;
DRAM[7680] = 8'b01100100;
DRAM[7681] = 8'b01100110;
DRAM[7682] = 8'b01100010;
DRAM[7683] = 8'b01100011;
DRAM[7684] = 8'b01100000;
DRAM[7685] = 8'b01011001;
DRAM[7686] = 8'b01100010;
DRAM[7687] = 8'b10000111;
DRAM[7688] = 8'b10011011;
DRAM[7689] = 8'b10100111;
DRAM[7690] = 8'b10101101;
DRAM[7691] = 8'b10101111;
DRAM[7692] = 8'b10101111;
DRAM[7693] = 8'b10101010;
DRAM[7694] = 8'b10011000;
DRAM[7695] = 8'b01111000;
DRAM[7696] = 8'b01010000;
DRAM[7697] = 8'b01001100;
DRAM[7698] = 8'b01011000;
DRAM[7699] = 8'b01100001;
DRAM[7700] = 8'b01100100;
DRAM[7701] = 8'b01100110;
DRAM[7702] = 8'b01100111;
DRAM[7703] = 8'b01100101;
DRAM[7704] = 8'b01100111;
DRAM[7705] = 8'b01100110;
DRAM[7706] = 8'b01101011;
DRAM[7707] = 8'b01101110;
DRAM[7708] = 8'b01110100;
DRAM[7709] = 8'b01111000;
DRAM[7710] = 8'b01111000;
DRAM[7711] = 8'b01111001;
DRAM[7712] = 8'b01111101;
DRAM[7713] = 8'b10000110;
DRAM[7714] = 8'b10010010;
DRAM[7715] = 8'b10011010;
DRAM[7716] = 8'b01111101;
DRAM[7717] = 8'b10000010;
DRAM[7718] = 8'b01111001;
DRAM[7719] = 8'b01011000;
DRAM[7720] = 8'b00111010;
DRAM[7721] = 8'b01010011;
DRAM[7722] = 8'b00100110;
DRAM[7723] = 8'b01110010;
DRAM[7724] = 8'b00101000;
DRAM[7725] = 8'b00110001;
DRAM[7726] = 8'b01010110;
DRAM[7727] = 8'b01001110;
DRAM[7728] = 8'b00110100;
DRAM[7729] = 8'b00101000;
DRAM[7730] = 8'b00110000;
DRAM[7731] = 8'b00111011;
DRAM[7732] = 8'b00101111;
DRAM[7733] = 8'b01001110;
DRAM[7734] = 8'b01000100;
DRAM[7735] = 8'b00101110;
DRAM[7736] = 8'b00110101;
DRAM[7737] = 8'b10000110;
DRAM[7738] = 8'b01110110;
DRAM[7739] = 8'b10101110;
DRAM[7740] = 8'b10101010;
DRAM[7741] = 8'b10100010;
DRAM[7742] = 8'b10101001;
DRAM[7743] = 8'b10111110;
DRAM[7744] = 8'b10111001;
DRAM[7745] = 8'b10110011;
DRAM[7746] = 8'b10011101;
DRAM[7747] = 8'b10000101;
DRAM[7748] = 8'b10010111;
DRAM[7749] = 8'b10100001;
DRAM[7750] = 8'b10100111;
DRAM[7751] = 8'b10101010;
DRAM[7752] = 8'b10110001;
DRAM[7753] = 8'b10110010;
DRAM[7754] = 8'b10110000;
DRAM[7755] = 8'b10110101;
DRAM[7756] = 8'b10111100;
DRAM[7757] = 8'b11000010;
DRAM[7758] = 8'b11000100;
DRAM[7759] = 8'b11000100;
DRAM[7760] = 8'b11000111;
DRAM[7761] = 8'b11001010;
DRAM[7762] = 8'b11001110;
DRAM[7763] = 8'b11010010;
DRAM[7764] = 8'b11010000;
DRAM[7765] = 8'b11000000;
DRAM[7766] = 8'b01111110;
DRAM[7767] = 8'b01000000;
DRAM[7768] = 8'b00100111;
DRAM[7769] = 8'b00101100;
DRAM[7770] = 8'b01000000;
DRAM[7771] = 8'b10110100;
DRAM[7772] = 8'b01010111;
DRAM[7773] = 8'b00111111;
DRAM[7774] = 8'b00111101;
DRAM[7775] = 8'b00111011;
DRAM[7776] = 8'b00111100;
DRAM[7777] = 8'b00111101;
DRAM[7778] = 8'b00110000;
DRAM[7779] = 8'b00110111;
DRAM[7780] = 8'b00110101;
DRAM[7781] = 8'b00101011;
DRAM[7782] = 8'b01001100;
DRAM[7783] = 8'b10000100;
DRAM[7784] = 8'b10000100;
DRAM[7785] = 8'b10001110;
DRAM[7786] = 8'b10100001;
DRAM[7787] = 8'b10100011;
DRAM[7788] = 8'b10100010;
DRAM[7789] = 8'b10100000;
DRAM[7790] = 8'b10100000;
DRAM[7791] = 8'b10100011;
DRAM[7792] = 8'b10100100;
DRAM[7793] = 8'b10100101;
DRAM[7794] = 8'b10100000;
DRAM[7795] = 8'b10011110;
DRAM[7796] = 8'b10011100;
DRAM[7797] = 8'b10010111;
DRAM[7798] = 8'b10010101;
DRAM[7799] = 8'b10010001;
DRAM[7800] = 8'b10001111;
DRAM[7801] = 8'b10010000;
DRAM[7802] = 8'b10010000;
DRAM[7803] = 8'b10001111;
DRAM[7804] = 8'b10001111;
DRAM[7805] = 8'b10001111;
DRAM[7806] = 8'b10010000;
DRAM[7807] = 8'b10010101;
DRAM[7808] = 8'b01100011;
DRAM[7809] = 8'b01100011;
DRAM[7810] = 8'b01100011;
DRAM[7811] = 8'b01100010;
DRAM[7812] = 8'b01100010;
DRAM[7813] = 8'b01011100;
DRAM[7814] = 8'b01100010;
DRAM[7815] = 8'b10000100;
DRAM[7816] = 8'b10011011;
DRAM[7817] = 8'b10100111;
DRAM[7818] = 8'b10110000;
DRAM[7819] = 8'b10110001;
DRAM[7820] = 8'b10101111;
DRAM[7821] = 8'b10101000;
DRAM[7822] = 8'b10010111;
DRAM[7823] = 8'b01110110;
DRAM[7824] = 8'b01010010;
DRAM[7825] = 8'b01001110;
DRAM[7826] = 8'b01011010;
DRAM[7827] = 8'b01011101;
DRAM[7828] = 8'b01100101;
DRAM[7829] = 8'b01100110;
DRAM[7830] = 8'b01100100;
DRAM[7831] = 8'b01100110;
DRAM[7832] = 8'b01100011;
DRAM[7833] = 8'b01100111;
DRAM[7834] = 8'b01101011;
DRAM[7835] = 8'b01110010;
DRAM[7836] = 8'b01110110;
DRAM[7837] = 8'b01111000;
DRAM[7838] = 8'b01111000;
DRAM[7839] = 8'b10101100;
DRAM[7840] = 8'b01110110;
DRAM[7841] = 8'b00101101;
DRAM[7842] = 8'b00100110;
DRAM[7843] = 8'b01101000;
DRAM[7844] = 8'b10101101;
DRAM[7845] = 8'b01101110;
DRAM[7846] = 8'b01100000;
DRAM[7847] = 8'b00111011;
DRAM[7848] = 8'b01100010;
DRAM[7849] = 8'b00101101;
DRAM[7850] = 8'b01000000;
DRAM[7851] = 8'b01001100;
DRAM[7852] = 8'b00101111;
DRAM[7853] = 8'b00110010;
DRAM[7854] = 8'b00110100;
DRAM[7855] = 8'b00110111;
DRAM[7856] = 8'b00101100;
DRAM[7857] = 8'b00110001;
DRAM[7858] = 8'b00110110;
DRAM[7859] = 8'b00111101;
DRAM[7860] = 8'b01001010;
DRAM[7861] = 8'b01001010;
DRAM[7862] = 8'b01000011;
DRAM[7863] = 8'b00100100;
DRAM[7864] = 8'b01110000;
DRAM[7865] = 8'b01101110;
DRAM[7866] = 8'b10101101;
DRAM[7867] = 8'b10101101;
DRAM[7868] = 8'b10111010;
DRAM[7869] = 8'b10011011;
DRAM[7870] = 8'b10101010;
DRAM[7871] = 8'b11000001;
DRAM[7872] = 8'b11000100;
DRAM[7873] = 8'b10000101;
DRAM[7874] = 8'b01100000;
DRAM[7875] = 8'b01101000;
DRAM[7876] = 8'b01101000;
DRAM[7877] = 8'b01101001;
DRAM[7878] = 8'b10000000;
DRAM[7879] = 8'b10011101;
DRAM[7880] = 8'b10101110;
DRAM[7881] = 8'b10110100;
DRAM[7882] = 8'b10110000;
DRAM[7883] = 8'b10101110;
DRAM[7884] = 8'b10110110;
DRAM[7885] = 8'b10111111;
DRAM[7886] = 8'b11000001;
DRAM[7887] = 8'b10111111;
DRAM[7888] = 8'b11000011;
DRAM[7889] = 8'b11001000;
DRAM[7890] = 8'b11001010;
DRAM[7891] = 8'b11001110;
DRAM[7892] = 8'b11000011;
DRAM[7893] = 8'b10011110;
DRAM[7894] = 8'b01011110;
DRAM[7895] = 8'b00110101;
DRAM[7896] = 8'b00100111;
DRAM[7897] = 8'b00100111;
DRAM[7898] = 8'b00110110;
DRAM[7899] = 8'b10100101;
DRAM[7900] = 8'b01101011;
DRAM[7901] = 8'b00111011;
DRAM[7902] = 8'b00111101;
DRAM[7903] = 8'b00111011;
DRAM[7904] = 8'b01000011;
DRAM[7905] = 8'b00111001;
DRAM[7906] = 8'b00110000;
DRAM[7907] = 8'b00110011;
DRAM[7908] = 8'b00110100;
DRAM[7909] = 8'b00101101;
DRAM[7910] = 8'b01100010;
DRAM[7911] = 8'b10001010;
DRAM[7912] = 8'b10000011;
DRAM[7913] = 8'b10011011;
DRAM[7914] = 8'b10100000;
DRAM[7915] = 8'b10100000;
DRAM[7916] = 8'b10011111;
DRAM[7917] = 8'b10011110;
DRAM[7918] = 8'b10100000;
DRAM[7919] = 8'b10100000;
DRAM[7920] = 8'b10011110;
DRAM[7921] = 8'b10100010;
DRAM[7922] = 8'b10100001;
DRAM[7923] = 8'b10011110;
DRAM[7924] = 8'b10011011;
DRAM[7925] = 8'b10011100;
DRAM[7926] = 8'b10011001;
DRAM[7927] = 8'b10010111;
DRAM[7928] = 8'b10010110;
DRAM[7929] = 8'b10010110;
DRAM[7930] = 8'b10010010;
DRAM[7931] = 8'b10001110;
DRAM[7932] = 8'b10001101;
DRAM[7933] = 8'b10001101;
DRAM[7934] = 8'b10001100;
DRAM[7935] = 8'b10001010;
DRAM[7936] = 8'b01100111;
DRAM[7937] = 8'b01100100;
DRAM[7938] = 8'b01100110;
DRAM[7939] = 8'b01100011;
DRAM[7940] = 8'b01100100;
DRAM[7941] = 8'b01011101;
DRAM[7942] = 8'b01100010;
DRAM[7943] = 8'b10000110;
DRAM[7944] = 8'b10011010;
DRAM[7945] = 8'b10101011;
DRAM[7946] = 8'b10101111;
DRAM[7947] = 8'b10110000;
DRAM[7948] = 8'b10110010;
DRAM[7949] = 8'b10101011;
DRAM[7950] = 8'b10011000;
DRAM[7951] = 8'b01111000;
DRAM[7952] = 8'b01001111;
DRAM[7953] = 8'b01010001;
DRAM[7954] = 8'b01011001;
DRAM[7955] = 8'b01011111;
DRAM[7956] = 8'b01100100;
DRAM[7957] = 8'b01101000;
DRAM[7958] = 8'b01100101;
DRAM[7959] = 8'b01100101;
DRAM[7960] = 8'b01100101;
DRAM[7961] = 8'b01100110;
DRAM[7962] = 8'b01101010;
DRAM[7963] = 8'b01101111;
DRAM[7964] = 8'b01110011;
DRAM[7965] = 8'b01110110;
DRAM[7966] = 8'b10000100;
DRAM[7967] = 8'b10010110;
DRAM[7968] = 8'b01101110;
DRAM[7969] = 8'b00110011;
DRAM[7970] = 8'b00100100;
DRAM[7971] = 8'b10001111;
DRAM[7972] = 8'b01101111;
DRAM[7973] = 8'b01010011;
DRAM[7974] = 8'b01001011;
DRAM[7975] = 8'b01001110;
DRAM[7976] = 8'b01001001;
DRAM[7977] = 8'b00101111;
DRAM[7978] = 8'b01010100;
DRAM[7979] = 8'b01011100;
DRAM[7980] = 8'b00100110;
DRAM[7981] = 8'b01000010;
DRAM[7982] = 8'b01000000;
DRAM[7983] = 8'b01000110;
DRAM[7984] = 8'b00110101;
DRAM[7985] = 8'b00101001;
DRAM[7986] = 8'b00101000;
DRAM[7987] = 8'b01001001;
DRAM[7988] = 8'b01010100;
DRAM[7989] = 8'b00111110;
DRAM[7990] = 8'b00101110;
DRAM[7991] = 8'b01011101;
DRAM[7992] = 8'b01111001;
DRAM[7993] = 8'b10101000;
DRAM[7994] = 8'b10101011;
DRAM[7995] = 8'b10111100;
DRAM[7996] = 8'b10110110;
DRAM[7997] = 8'b10011100;
DRAM[7998] = 8'b10111010;
DRAM[7999] = 8'b11000011;
DRAM[8000] = 8'b10001011;
DRAM[8001] = 8'b10001101;
DRAM[8002] = 8'b10010101;
DRAM[8003] = 8'b10011001;
DRAM[8004] = 8'b10001001;
DRAM[8005] = 8'b01100100;
DRAM[8006] = 8'b01001110;
DRAM[8007] = 8'b01001010;
DRAM[8008] = 8'b01101110;
DRAM[8009] = 8'b10100000;
DRAM[8010] = 8'b10101100;
DRAM[8011] = 8'b10101010;
DRAM[8012] = 8'b10110000;
DRAM[8013] = 8'b10111110;
DRAM[8014] = 8'b11000001;
DRAM[8015] = 8'b10111110;
DRAM[8016] = 8'b11000001;
DRAM[8017] = 8'b11000001;
DRAM[8018] = 8'b10110110;
DRAM[8019] = 8'b10001100;
DRAM[8020] = 8'b01101100;
DRAM[8021] = 8'b01100011;
DRAM[8022] = 8'b01011110;
DRAM[8023] = 8'b01001100;
DRAM[8024] = 8'b00101111;
DRAM[8025] = 8'b00101010;
DRAM[8026] = 8'b00111001;
DRAM[8027] = 8'b10011100;
DRAM[8028] = 8'b01111110;
DRAM[8029] = 8'b00111010;
DRAM[8030] = 8'b00111011;
DRAM[8031] = 8'b00111111;
DRAM[8032] = 8'b00111110;
DRAM[8033] = 8'b00110100;
DRAM[8034] = 8'b00110010;
DRAM[8035] = 8'b00110100;
DRAM[8036] = 8'b00111001;
DRAM[8037] = 8'b00110011;
DRAM[8038] = 8'b01110110;
DRAM[8039] = 8'b10000111;
DRAM[8040] = 8'b10001000;
DRAM[8041] = 8'b10011111;
DRAM[8042] = 8'b10100001;
DRAM[8043] = 8'b10011110;
DRAM[8044] = 8'b10011100;
DRAM[8045] = 8'b10011110;
DRAM[8046] = 8'b10011011;
DRAM[8047] = 8'b10011100;
DRAM[8048] = 8'b10011011;
DRAM[8049] = 8'b10011011;
DRAM[8050] = 8'b10011101;
DRAM[8051] = 8'b10011011;
DRAM[8052] = 8'b10011011;
DRAM[8053] = 8'b10011010;
DRAM[8054] = 8'b10011001;
DRAM[8055] = 8'b10011010;
DRAM[8056] = 8'b10011100;
DRAM[8057] = 8'b10011010;
DRAM[8058] = 8'b10011000;
DRAM[8059] = 8'b10010010;
DRAM[8060] = 8'b10001111;
DRAM[8061] = 8'b10001101;
DRAM[8062] = 8'b10001000;
DRAM[8063] = 8'b10000100;
DRAM[8064] = 8'b01100100;
DRAM[8065] = 8'b01100111;
DRAM[8066] = 8'b01101011;
DRAM[8067] = 8'b01100111;
DRAM[8068] = 8'b01100010;
DRAM[8069] = 8'b01011011;
DRAM[8070] = 8'b01100001;
DRAM[8071] = 8'b10000101;
DRAM[8072] = 8'b10011001;
DRAM[8073] = 8'b10101001;
DRAM[8074] = 8'b10101110;
DRAM[8075] = 8'b10110000;
DRAM[8076] = 8'b10110001;
DRAM[8077] = 8'b10101100;
DRAM[8078] = 8'b10011001;
DRAM[8079] = 8'b01111011;
DRAM[8080] = 8'b01010011;
DRAM[8081] = 8'b01010001;
DRAM[8082] = 8'b01011001;
DRAM[8083] = 8'b01100000;
DRAM[8084] = 8'b01100111;
DRAM[8085] = 8'b01100101;
DRAM[8086] = 8'b01100101;
DRAM[8087] = 8'b01100100;
DRAM[8088] = 8'b01100010;
DRAM[8089] = 8'b01100110;
DRAM[8090] = 8'b01100110;
DRAM[8091] = 8'b01101001;
DRAM[8092] = 8'b01110000;
DRAM[8093] = 8'b10000110;
DRAM[8094] = 8'b10011100;
DRAM[8095] = 8'b10010010;
DRAM[8096] = 8'b10011001;
DRAM[8097] = 8'b01111000;
DRAM[8098] = 8'b01010110;
DRAM[8099] = 8'b10000000;
DRAM[8100] = 8'b01100001;
DRAM[8101] = 8'b00111101;
DRAM[8102] = 8'b00111111;
DRAM[8103] = 8'b01100001;
DRAM[8104] = 8'b00111111;
DRAM[8105] = 8'b01011110;
DRAM[8106] = 8'b00101111;
DRAM[8107] = 8'b01100000;
DRAM[8108] = 8'b00101010;
DRAM[8109] = 8'b00111100;
DRAM[8110] = 8'b00101000;
DRAM[8111] = 8'b00111101;
DRAM[8112] = 8'b01001011;
DRAM[8113] = 8'b00101000;
DRAM[8114] = 8'b00101110;
DRAM[8115] = 8'b00101011;
DRAM[8116] = 8'b00111111;
DRAM[8117] = 8'b00110010;
DRAM[8118] = 8'b00101110;
DRAM[8119] = 8'b10000111;
DRAM[8120] = 8'b10011000;
DRAM[8121] = 8'b10101011;
DRAM[8122] = 8'b10110111;
DRAM[8123] = 8'b11000101;
DRAM[8124] = 8'b10101010;
DRAM[8125] = 8'b10101111;
DRAM[8126] = 8'b10110010;
DRAM[8127] = 8'b01110101;
DRAM[8128] = 8'b01101110;
DRAM[8129] = 8'b01110011;
DRAM[8130] = 8'b01110100;
DRAM[8131] = 8'b01100000;
DRAM[8132] = 8'b01111110;
DRAM[8133] = 8'b01101100;
DRAM[8134] = 8'b01110000;
DRAM[8135] = 8'b01100100;
DRAM[8136] = 8'b01100010;
DRAM[8137] = 8'b01111010;
DRAM[8138] = 8'b10011110;
DRAM[8139] = 8'b10100011;
DRAM[8140] = 8'b10101010;
DRAM[8141] = 8'b10111100;
DRAM[8142] = 8'b11000010;
DRAM[8143] = 8'b10111101;
DRAM[8144] = 8'b10111011;
DRAM[8145] = 8'b10100100;
DRAM[8146] = 8'b01110100;
DRAM[8147] = 8'b01101010;
DRAM[8148] = 8'b01101000;
DRAM[8149] = 8'b01101000;
DRAM[8150] = 8'b01100010;
DRAM[8151] = 8'b01010000;
DRAM[8152] = 8'b00111010;
DRAM[8153] = 8'b00101011;
DRAM[8154] = 8'b00111111;
DRAM[8155] = 8'b10001111;
DRAM[8156] = 8'b10000000;
DRAM[8157] = 8'b00111110;
DRAM[8158] = 8'b01000100;
DRAM[8159] = 8'b00111100;
DRAM[8160] = 8'b01000001;
DRAM[8161] = 8'b00110000;
DRAM[8162] = 8'b00111000;
DRAM[8163] = 8'b00110100;
DRAM[8164] = 8'b00110101;
DRAM[8165] = 8'b01001000;
DRAM[8166] = 8'b10000110;
DRAM[8167] = 8'b10000101;
DRAM[8168] = 8'b10010001;
DRAM[8169] = 8'b10100000;
DRAM[8170] = 8'b10011110;
DRAM[8171] = 8'b10011101;
DRAM[8172] = 8'b10011011;
DRAM[8173] = 8'b10011110;
DRAM[8174] = 8'b10011110;
DRAM[8175] = 8'b10011011;
DRAM[8176] = 8'b10011101;
DRAM[8177] = 8'b10011110;
DRAM[8178] = 8'b10011111;
DRAM[8179] = 8'b10011100;
DRAM[8180] = 8'b10011100;
DRAM[8181] = 8'b10011000;
DRAM[8182] = 8'b10011011;
DRAM[8183] = 8'b10011010;
DRAM[8184] = 8'b10011100;
DRAM[8185] = 8'b10011100;
DRAM[8186] = 8'b10011010;
DRAM[8187] = 8'b10010110;
DRAM[8188] = 8'b10010111;
DRAM[8189] = 8'b10001111;
DRAM[8190] = 8'b10000111;
DRAM[8191] = 8'b10000101;
DRAM[8192] = 8'b01100110;
DRAM[8193] = 8'b01100110;
DRAM[8194] = 8'b01100100;
DRAM[8195] = 8'b01100100;
DRAM[8196] = 8'b01011111;
DRAM[8197] = 8'b01011001;
DRAM[8198] = 8'b01011110;
DRAM[8199] = 8'b10000100;
DRAM[8200] = 8'b10011010;
DRAM[8201] = 8'b10101010;
DRAM[8202] = 8'b10110001;
DRAM[8203] = 8'b10110000;
DRAM[8204] = 8'b10101111;
DRAM[8205] = 8'b10101010;
DRAM[8206] = 8'b10011010;
DRAM[8207] = 8'b01111001;
DRAM[8208] = 8'b01010000;
DRAM[8209] = 8'b01001100;
DRAM[8210] = 8'b01010100;
DRAM[8211] = 8'b01100000;
DRAM[8212] = 8'b01100101;
DRAM[8213] = 8'b01100110;
DRAM[8214] = 8'b01100100;
DRAM[8215] = 8'b01100100;
DRAM[8216] = 8'b01011111;
DRAM[8217] = 8'b01100000;
DRAM[8218] = 8'b01100001;
DRAM[8219] = 8'b01111101;
DRAM[8220] = 8'b10010110;
DRAM[8221] = 8'b10010010;
DRAM[8222] = 8'b10011010;
DRAM[8223] = 8'b10011011;
DRAM[8224] = 8'b10011010;
DRAM[8225] = 8'b01111101;
DRAM[8226] = 8'b01101010;
DRAM[8227] = 8'b00101110;
DRAM[8228] = 8'b00101101;
DRAM[8229] = 8'b01010010;
DRAM[8230] = 8'b01100011;
DRAM[8231] = 8'b01010000;
DRAM[8232] = 8'b01010001;
DRAM[8233] = 8'b01100100;
DRAM[8234] = 8'b00100011;
DRAM[8235] = 8'b00110000;
DRAM[8236] = 8'b00110110;
DRAM[8237] = 8'b01001011;
DRAM[8238] = 8'b00101001;
DRAM[8239] = 8'b00101001;
DRAM[8240] = 8'b01011000;
DRAM[8241] = 8'b00111100;
DRAM[8242] = 8'b00101010;
DRAM[8243] = 8'b00101101;
DRAM[8244] = 8'b00101001;
DRAM[8245] = 8'b00011111;
DRAM[8246] = 8'b01110001;
DRAM[8247] = 8'b01111010;
DRAM[8248] = 8'b10110010;
DRAM[8249] = 8'b10110000;
DRAM[8250] = 8'b11000110;
DRAM[8251] = 8'b11000000;
DRAM[8252] = 8'b10110110;
DRAM[8253] = 8'b10101011;
DRAM[8254] = 8'b01001000;
DRAM[8255] = 8'b01001010;
DRAM[8256] = 8'b00111111;
DRAM[8257] = 8'b00111001;
DRAM[8258] = 8'b00110011;
DRAM[8259] = 8'b00110000;
DRAM[8260] = 8'b00110110;
DRAM[8261] = 8'b00101100;
DRAM[8262] = 8'b01000100;
DRAM[8263] = 8'b10000111;
DRAM[8264] = 8'b01111110;
DRAM[8265] = 8'b01111110;
DRAM[8266] = 8'b10001110;
DRAM[8267] = 8'b10011011;
DRAM[8268] = 8'b10100101;
DRAM[8269] = 8'b10111101;
DRAM[8270] = 8'b11000011;
DRAM[8271] = 8'b11000101;
DRAM[8272] = 8'b10110101;
DRAM[8273] = 8'b01110101;
DRAM[8274] = 8'b01001011;
DRAM[8275] = 8'b00110100;
DRAM[8276] = 8'b00110000;
DRAM[8277] = 8'b00110110;
DRAM[8278] = 8'b00111010;
DRAM[8279] = 8'b01000000;
DRAM[8280] = 8'b00110100;
DRAM[8281] = 8'b00101000;
DRAM[8282] = 8'b00111111;
DRAM[8283] = 8'b01111011;
DRAM[8284] = 8'b10001010;
DRAM[8285] = 8'b01000110;
DRAM[8286] = 8'b01000001;
DRAM[8287] = 8'b00111100;
DRAM[8288] = 8'b00110011;
DRAM[8289] = 8'b00101111;
DRAM[8290] = 8'b00110011;
DRAM[8291] = 8'b00110101;
DRAM[8292] = 8'b00101010;
DRAM[8293] = 8'b01010110;
DRAM[8294] = 8'b10001101;
DRAM[8295] = 8'b10000100;
DRAM[8296] = 8'b10011000;
DRAM[8297] = 8'b10100000;
DRAM[8298] = 8'b10011111;
DRAM[8299] = 8'b10011010;
DRAM[8300] = 8'b10011010;
DRAM[8301] = 8'b10011100;
DRAM[8302] = 8'b10011010;
DRAM[8303] = 8'b10011101;
DRAM[8304] = 8'b10011100;
DRAM[8305] = 8'b10011011;
DRAM[8306] = 8'b10011100;
DRAM[8307] = 8'b10011101;
DRAM[8308] = 8'b10011001;
DRAM[8309] = 8'b10011001;
DRAM[8310] = 8'b10011010;
DRAM[8311] = 8'b10011010;
DRAM[8312] = 8'b10011001;
DRAM[8313] = 8'b10011100;
DRAM[8314] = 8'b10010111;
DRAM[8315] = 8'b10010011;
DRAM[8316] = 8'b10010000;
DRAM[8317] = 8'b10010000;
DRAM[8318] = 8'b10001010;
DRAM[8319] = 8'b10001000;
DRAM[8320] = 8'b01011111;
DRAM[8321] = 8'b01100000;
DRAM[8322] = 8'b01100000;
DRAM[8323] = 8'b01011110;
DRAM[8324] = 8'b01011001;
DRAM[8325] = 8'b01001111;
DRAM[8326] = 8'b01011010;
DRAM[8327] = 8'b10000000;
DRAM[8328] = 8'b10011000;
DRAM[8329] = 8'b10101000;
DRAM[8330] = 8'b10101111;
DRAM[8331] = 8'b10110010;
DRAM[8332] = 8'b10110000;
DRAM[8333] = 8'b10101001;
DRAM[8334] = 8'b10010111;
DRAM[8335] = 8'b01111011;
DRAM[8336] = 8'b01001110;
DRAM[8337] = 8'b01001000;
DRAM[8338] = 8'b01010110;
DRAM[8339] = 8'b01011101;
DRAM[8340] = 8'b01011111;
DRAM[8341] = 8'b01100011;
DRAM[8342] = 8'b01100100;
DRAM[8343] = 8'b01011110;
DRAM[8344] = 8'b01011101;
DRAM[8345] = 8'b01010111;
DRAM[8346] = 8'b10000010;
DRAM[8347] = 8'b11000100;
DRAM[8348] = 8'b10011101;
DRAM[8349] = 8'b10010001;
DRAM[8350] = 8'b10011000;
DRAM[8351] = 8'b10001010;
DRAM[8352] = 8'b01111100;
DRAM[8353] = 8'b01000100;
DRAM[8354] = 8'b00110110;
DRAM[8355] = 8'b00100100;
DRAM[8356] = 8'b01101100;
DRAM[8357] = 8'b01000101;
DRAM[8358] = 8'b01010111;
DRAM[8359] = 8'b01000101;
DRAM[8360] = 8'b01010000;
DRAM[8361] = 8'b01111000;
DRAM[8362] = 8'b00100100;
DRAM[8363] = 8'b00111001;
DRAM[8364] = 8'b00111000;
DRAM[8365] = 8'b01011101;
DRAM[8366] = 8'b00101001;
DRAM[8367] = 8'b00101000;
DRAM[8368] = 8'b00101010;
DRAM[8369] = 8'b01100110;
DRAM[8370] = 8'b01001110;
DRAM[8371] = 8'b00100111;
DRAM[8372] = 8'b00100100;
DRAM[8373] = 8'b01000101;
DRAM[8374] = 8'b01111000;
DRAM[8375] = 8'b10110010;
DRAM[8376] = 8'b10101010;
DRAM[8377] = 8'b10110100;
DRAM[8378] = 8'b11000110;
DRAM[8379] = 8'b11000000;
DRAM[8380] = 8'b10101011;
DRAM[8381] = 8'b01000110;
DRAM[8382] = 8'b00111011;
DRAM[8383] = 8'b00110001;
DRAM[8384] = 8'b00110011;
DRAM[8385] = 8'b00110010;
DRAM[8386] = 8'b00110101;
DRAM[8387] = 8'b01001101;
DRAM[8388] = 8'b10010110;
DRAM[8389] = 8'b01000001;
DRAM[8390] = 8'b00101000;
DRAM[8391] = 8'b01001001;
DRAM[8392] = 8'b10000101;
DRAM[8393] = 8'b01111110;
DRAM[8394] = 8'b10001100;
DRAM[8395] = 8'b10010110;
DRAM[8396] = 8'b10100101;
DRAM[8397] = 8'b11000001;
DRAM[8398] = 8'b11001111;
DRAM[8399] = 8'b11000110;
DRAM[8400] = 8'b01010001;
DRAM[8401] = 8'b00110001;
DRAM[8402] = 8'b00111111;
DRAM[8403] = 8'b01100111;
DRAM[8404] = 8'b01011101;
DRAM[8405] = 8'b00101110;
DRAM[8406] = 8'b00111000;
DRAM[8407] = 8'b00111000;
DRAM[8408] = 8'b00101110;
DRAM[8409] = 8'b00101010;
DRAM[8410] = 8'b00111000;
DRAM[8411] = 8'b01101101;
DRAM[8412] = 8'b01111111;
DRAM[8413] = 8'b01010010;
DRAM[8414] = 8'b01001000;
DRAM[8415] = 8'b00111100;
DRAM[8416] = 8'b00110001;
DRAM[8417] = 8'b00110001;
DRAM[8418] = 8'b00110000;
DRAM[8419] = 8'b00110010;
DRAM[8420] = 8'b00101110;
DRAM[8421] = 8'b01110100;
DRAM[8422] = 8'b10001100;
DRAM[8423] = 8'b10001110;
DRAM[8424] = 8'b10100001;
DRAM[8425] = 8'b10011110;
DRAM[8426] = 8'b10011011;
DRAM[8427] = 8'b10011001;
DRAM[8428] = 8'b10011001;
DRAM[8429] = 8'b10011010;
DRAM[8430] = 8'b10011011;
DRAM[8431] = 8'b10011011;
DRAM[8432] = 8'b10011001;
DRAM[8433] = 8'b10011100;
DRAM[8434] = 8'b10011001;
DRAM[8435] = 8'b10011001;
DRAM[8436] = 8'b10011011;
DRAM[8437] = 8'b10011010;
DRAM[8438] = 8'b10011000;
DRAM[8439] = 8'b10010100;
DRAM[8440] = 8'b10010111;
DRAM[8441] = 8'b10010101;
DRAM[8442] = 8'b10001111;
DRAM[8443] = 8'b10001110;
DRAM[8444] = 8'b10001010;
DRAM[8445] = 8'b10001011;
DRAM[8446] = 8'b10001000;
DRAM[8447] = 8'b10000111;
DRAM[8448] = 8'b01100100;
DRAM[8449] = 8'b01100000;
DRAM[8450] = 8'b01100000;
DRAM[8451] = 8'b01011101;
DRAM[8452] = 8'b01010110;
DRAM[8453] = 8'b01001110;
DRAM[8454] = 8'b01010100;
DRAM[8455] = 8'b01111111;
DRAM[8456] = 8'b10011001;
DRAM[8457] = 8'b10101100;
DRAM[8458] = 8'b10110001;
DRAM[8459] = 8'b10110001;
DRAM[8460] = 8'b10110010;
DRAM[8461] = 8'b10101011;
DRAM[8462] = 8'b10011000;
DRAM[8463] = 8'b01111010;
DRAM[8464] = 8'b01001110;
DRAM[8465] = 8'b01001110;
DRAM[8466] = 8'b01011001;
DRAM[8467] = 8'b01100011;
DRAM[8468] = 8'b01100011;
DRAM[8469] = 8'b01100010;
DRAM[8470] = 8'b01100011;
DRAM[8471] = 8'b01100100;
DRAM[8472] = 8'b01011110;
DRAM[8473] = 8'b01011000;
DRAM[8474] = 8'b01111100;
DRAM[8475] = 8'b10110011;
DRAM[8476] = 8'b10011011;
DRAM[8477] = 8'b10010000;
DRAM[8478] = 8'b10010111;
DRAM[8479] = 8'b10000001;
DRAM[8480] = 8'b01101111;
DRAM[8481] = 8'b00101111;
DRAM[8482] = 8'b00110010;
DRAM[8483] = 8'b01010010;
DRAM[8484] = 8'b00110000;
DRAM[8485] = 8'b01001010;
DRAM[8486] = 8'b00101111;
DRAM[8487] = 8'b01000100;
DRAM[8488] = 8'b01100011;
DRAM[8489] = 8'b01011001;
DRAM[8490] = 8'b00101101;
DRAM[8491] = 8'b00101101;
DRAM[8492] = 8'b00101110;
DRAM[8493] = 8'b01001010;
DRAM[8494] = 8'b00111110;
DRAM[8495] = 8'b00101010;
DRAM[8496] = 8'b00101101;
DRAM[8497] = 8'b00110000;
DRAM[8498] = 8'b00110010;
DRAM[8499] = 8'b00110011;
DRAM[8500] = 8'b00101111;
DRAM[8501] = 8'b01111100;
DRAM[8502] = 8'b10001101;
DRAM[8503] = 8'b10110001;
DRAM[8504] = 8'b10110011;
DRAM[8505] = 8'b11000000;
DRAM[8506] = 8'b11001001;
DRAM[8507] = 8'b10111010;
DRAM[8508] = 8'b01011010;
DRAM[8509] = 8'b01001011;
DRAM[8510] = 8'b00110000;
DRAM[8511] = 8'b00111000;
DRAM[8512] = 8'b01010000;
DRAM[8513] = 8'b01001110;
DRAM[8514] = 8'b00111011;
DRAM[8515] = 8'b00111110;
DRAM[8516] = 8'b11001101;
DRAM[8517] = 8'b10110110;
DRAM[8518] = 8'b01010001;
DRAM[8519] = 8'b01100110;
DRAM[8520] = 8'b01110101;
DRAM[8521] = 8'b01111000;
DRAM[8522] = 8'b10000101;
DRAM[8523] = 8'b10010001;
DRAM[8524] = 8'b10100101;
DRAM[8525] = 8'b11000111;
DRAM[8526] = 8'b11010111;
DRAM[8527] = 8'b01111000;
DRAM[8528] = 8'b00111100;
DRAM[8529] = 8'b00110101;
DRAM[8530] = 8'b01000010;
DRAM[8531] = 8'b10001011;
DRAM[8532] = 8'b10010101;
DRAM[8533] = 8'b00111101;
DRAM[8534] = 8'b00101110;
DRAM[8535] = 8'b00110000;
DRAM[8536] = 8'b00101100;
DRAM[8537] = 8'b00110010;
DRAM[8538] = 8'b00111111;
DRAM[8539] = 8'b01101010;
DRAM[8540] = 8'b10001101;
DRAM[8541] = 8'b01001110;
DRAM[8542] = 8'b01010001;
DRAM[8543] = 8'b00111001;
DRAM[8544] = 8'b00110010;
DRAM[8545] = 8'b00101110;
DRAM[8546] = 8'b00110110;
DRAM[8547] = 8'b00101110;
DRAM[8548] = 8'b01000010;
DRAM[8549] = 8'b10000110;
DRAM[8550] = 8'b10001110;
DRAM[8551] = 8'b10010011;
DRAM[8552] = 8'b10100000;
DRAM[8553] = 8'b10011101;
DRAM[8554] = 8'b10011110;
DRAM[8555] = 8'b10011010;
DRAM[8556] = 8'b10011010;
DRAM[8557] = 8'b10011001;
DRAM[8558] = 8'b10011000;
DRAM[8559] = 8'b10011010;
DRAM[8560] = 8'b10011000;
DRAM[8561] = 8'b10011000;
DRAM[8562] = 8'b10011000;
DRAM[8563] = 8'b10011010;
DRAM[8564] = 8'b10011000;
DRAM[8565] = 8'b10011001;
DRAM[8566] = 8'b10010101;
DRAM[8567] = 8'b10010110;
DRAM[8568] = 8'b10010100;
DRAM[8569] = 8'b10010000;
DRAM[8570] = 8'b10001110;
DRAM[8571] = 8'b10001010;
DRAM[8572] = 8'b10000110;
DRAM[8573] = 8'b10000101;
DRAM[8574] = 8'b10000001;
DRAM[8575] = 8'b10000110;
DRAM[8576] = 8'b01100011;
DRAM[8577] = 8'b01100011;
DRAM[8578] = 8'b01100000;
DRAM[8579] = 8'b01011100;
DRAM[8580] = 8'b01011100;
DRAM[8581] = 8'b01001100;
DRAM[8582] = 8'b01010010;
DRAM[8583] = 8'b01111101;
DRAM[8584] = 8'b10011001;
DRAM[8585] = 8'b10101100;
DRAM[8586] = 8'b10110100;
DRAM[8587] = 8'b10110011;
DRAM[8588] = 8'b10110101;
DRAM[8589] = 8'b10101101;
DRAM[8590] = 8'b10011000;
DRAM[8591] = 8'b01111000;
DRAM[8592] = 8'b01010101;
DRAM[8593] = 8'b01010010;
DRAM[8594] = 8'b01011101;
DRAM[8595] = 8'b01100100;
DRAM[8596] = 8'b01101001;
DRAM[8597] = 8'b01100111;
DRAM[8598] = 8'b01101000;
DRAM[8599] = 8'b01101010;
DRAM[8600] = 8'b01011110;
DRAM[8601] = 8'b00111111;
DRAM[8602] = 8'b01000010;
DRAM[8603] = 8'b10000101;
DRAM[8604] = 8'b10101001;
DRAM[8605] = 8'b11001101;
DRAM[8606] = 8'b10001100;
DRAM[8607] = 8'b00110100;
DRAM[8608] = 8'b00101011;
DRAM[8609] = 8'b00101001;
DRAM[8610] = 8'b01010100;
DRAM[8611] = 8'b00111110;
DRAM[8612] = 8'b01000011;
DRAM[8613] = 8'b00111110;
DRAM[8614] = 8'b01000110;
DRAM[8615] = 8'b01101010;
DRAM[8616] = 8'b01011011;
DRAM[8617] = 8'b01100111;
DRAM[8618] = 8'b00101010;
DRAM[8619] = 8'b00110000;
DRAM[8620] = 8'b00110001;
DRAM[8621] = 8'b00101111;
DRAM[8622] = 8'b01001011;
DRAM[8623] = 8'b00110001;
DRAM[8624] = 8'b00101011;
DRAM[8625] = 8'b00110001;
DRAM[8626] = 8'b00100110;
DRAM[8627] = 8'b00101001;
DRAM[8628] = 8'b01010011;
DRAM[8629] = 8'b01100100;
DRAM[8630] = 8'b10100000;
DRAM[8631] = 8'b10100100;
DRAM[8632] = 8'b10111010;
DRAM[8633] = 8'b11000111;
DRAM[8634] = 8'b10111110;
DRAM[8635] = 8'b01111000;
DRAM[8636] = 8'b01111001;
DRAM[8637] = 8'b01110100;
DRAM[8638] = 8'b01010101;
DRAM[8639] = 8'b00111111;
DRAM[8640] = 8'b01110001;
DRAM[8641] = 8'b01010011;
DRAM[8642] = 8'b01001100;
DRAM[8643] = 8'b10010101;
DRAM[8644] = 8'b11001111;
DRAM[8645] = 8'b11000111;
DRAM[8646] = 8'b10000101;
DRAM[8647] = 8'b01110000;
DRAM[8648] = 8'b01101101;
DRAM[8649] = 8'b01110111;
DRAM[8650] = 8'b10000000;
DRAM[8651] = 8'b10001111;
DRAM[8652] = 8'b10101010;
DRAM[8653] = 8'b11010010;
DRAM[8654] = 8'b11001110;
DRAM[8655] = 8'b01101001;
DRAM[8656] = 8'b01101100;
DRAM[8657] = 8'b01011000;
DRAM[8658] = 8'b01001111;
DRAM[8659] = 8'b10010000;
DRAM[8660] = 8'b10011001;
DRAM[8661] = 8'b01000101;
DRAM[8662] = 8'b00101110;
DRAM[8663] = 8'b00101111;
DRAM[8664] = 8'b00101100;
DRAM[8665] = 8'b00101100;
DRAM[8666] = 8'b00111101;
DRAM[8667] = 8'b01110100;
DRAM[8668] = 8'b10100010;
DRAM[8669] = 8'b01001111;
DRAM[8670] = 8'b01010010;
DRAM[8671] = 8'b00111010;
DRAM[8672] = 8'b00101111;
DRAM[8673] = 8'b00110100;
DRAM[8674] = 8'b00110101;
DRAM[8675] = 8'b00101101;
DRAM[8676] = 8'b01010001;
DRAM[8677] = 8'b10001100;
DRAM[8678] = 8'b10001011;
DRAM[8679] = 8'b10011010;
DRAM[8680] = 8'b10011101;
DRAM[8681] = 8'b10011010;
DRAM[8682] = 8'b10011100;
DRAM[8683] = 8'b10010111;
DRAM[8684] = 8'b10010111;
DRAM[8685] = 8'b10011000;
DRAM[8686] = 8'b10011000;
DRAM[8687] = 8'b10011001;
DRAM[8688] = 8'b10011011;
DRAM[8689] = 8'b10011001;
DRAM[8690] = 8'b10011001;
DRAM[8691] = 8'b10010110;
DRAM[8692] = 8'b10011001;
DRAM[8693] = 8'b10010010;
DRAM[8694] = 8'b10010101;
DRAM[8695] = 8'b10010011;
DRAM[8696] = 8'b10010000;
DRAM[8697] = 8'b10001100;
DRAM[8698] = 8'b10000111;
DRAM[8699] = 8'b10000101;
DRAM[8700] = 8'b10000011;
DRAM[8701] = 8'b10000110;
DRAM[8702] = 8'b10010110;
DRAM[8703] = 8'b10100101;
DRAM[8704] = 8'b01100101;
DRAM[8705] = 8'b01100100;
DRAM[8706] = 8'b01100010;
DRAM[8707] = 8'b01011100;
DRAM[8708] = 8'b01011000;
DRAM[8709] = 8'b01001110;
DRAM[8710] = 8'b01001110;
DRAM[8711] = 8'b01111101;
DRAM[8712] = 8'b10011010;
DRAM[8713] = 8'b10101001;
DRAM[8714] = 8'b10110010;
DRAM[8715] = 8'b10110100;
DRAM[8716] = 8'b10110100;
DRAM[8717] = 8'b10101111;
DRAM[8718] = 8'b10011001;
DRAM[8719] = 8'b01111010;
DRAM[8720] = 8'b01011010;
DRAM[8721] = 8'b01011000;
DRAM[8722] = 8'b01100000;
DRAM[8723] = 8'b01100110;
DRAM[8724] = 8'b01101111;
DRAM[8725] = 8'b01101111;
DRAM[8726] = 8'b01100101;
DRAM[8727] = 8'b00110111;
DRAM[8728] = 8'b00110011;
DRAM[8729] = 8'b01110011;
DRAM[8730] = 8'b10010101;
DRAM[8731] = 8'b10110001;
DRAM[8732] = 8'b11001000;
DRAM[8733] = 8'b10010001;
DRAM[8734] = 8'b00110001;
DRAM[8735] = 8'b00111101;
DRAM[8736] = 8'b00111011;
DRAM[8737] = 8'b01101010;
DRAM[8738] = 8'b01010000;
DRAM[8739] = 8'b00101111;
DRAM[8740] = 8'b01001010;
DRAM[8741] = 8'b01010000;
DRAM[8742] = 8'b01010010;
DRAM[8743] = 8'b01101001;
DRAM[8744] = 8'b01101010;
DRAM[8745] = 8'b10000010;
DRAM[8746] = 8'b00111000;
DRAM[8747] = 8'b00111010;
DRAM[8748] = 8'b00101001;
DRAM[8749] = 8'b00101010;
DRAM[8750] = 8'b00110011;
DRAM[8751] = 8'b00110101;
DRAM[8752] = 8'b00110000;
DRAM[8753] = 8'b00101101;
DRAM[8754] = 8'b00100110;
DRAM[8755] = 8'b00101100;
DRAM[8756] = 8'b10000001;
DRAM[8757] = 8'b10100111;
DRAM[8758] = 8'b10100001;
DRAM[8759] = 8'b10110111;
DRAM[8760] = 8'b11000111;
DRAM[8761] = 8'b10111001;
DRAM[8762] = 8'b01110011;
DRAM[8763] = 8'b01111101;
DRAM[8764] = 8'b01111100;
DRAM[8765] = 8'b10010000;
DRAM[8766] = 8'b10000011;
DRAM[8767] = 8'b01101010;
DRAM[8768] = 8'b01101100;
DRAM[8769] = 8'b10000001;
DRAM[8770] = 8'b10010110;
DRAM[8771] = 8'b10110001;
DRAM[8772] = 8'b10111101;
DRAM[8773] = 8'b10110100;
DRAM[8774] = 8'b10010111;
DRAM[8775] = 8'b01111111;
DRAM[8776] = 8'b01111101;
DRAM[8777] = 8'b01111000;
DRAM[8778] = 8'b10000001;
DRAM[8779] = 8'b10001010;
DRAM[8780] = 8'b10101010;
DRAM[8781] = 8'b11011000;
DRAM[8782] = 8'b10111101;
DRAM[8783] = 8'b01110011;
DRAM[8784] = 8'b01111111;
DRAM[8785] = 8'b10000111;
DRAM[8786] = 8'b10011011;
DRAM[8787] = 8'b10100011;
DRAM[8788] = 8'b01111111;
DRAM[8789] = 8'b00111010;
DRAM[8790] = 8'b00111101;
DRAM[8791] = 8'b00110110;
DRAM[8792] = 8'b00110001;
DRAM[8793] = 8'b00110110;
DRAM[8794] = 8'b01000110;
DRAM[8795] = 8'b01101110;
DRAM[8796] = 8'b10100110;
DRAM[8797] = 8'b01010100;
DRAM[8798] = 8'b01010100;
DRAM[8799] = 8'b00110100;
DRAM[8800] = 8'b00110010;
DRAM[8801] = 8'b00110000;
DRAM[8802] = 8'b00110101;
DRAM[8803] = 8'b00110000;
DRAM[8804] = 8'b01101101;
DRAM[8805] = 8'b10001101;
DRAM[8806] = 8'b10001011;
DRAM[8807] = 8'b10011111;
DRAM[8808] = 8'b10011101;
DRAM[8809] = 8'b10011011;
DRAM[8810] = 8'b10011000;
DRAM[8811] = 8'b10011000;
DRAM[8812] = 8'b10010100;
DRAM[8813] = 8'b10011001;
DRAM[8814] = 8'b10100011;
DRAM[8815] = 8'b10011000;
DRAM[8816] = 8'b10011000;
DRAM[8817] = 8'b10011010;
DRAM[8818] = 8'b10010110;
DRAM[8819] = 8'b10010101;
DRAM[8820] = 8'b10010101;
DRAM[8821] = 8'b10010011;
DRAM[8822] = 8'b10001111;
DRAM[8823] = 8'b10001100;
DRAM[8824] = 8'b10001011;
DRAM[8825] = 8'b10001100;
DRAM[8826] = 8'b10000100;
DRAM[8827] = 8'b10001011;
DRAM[8828] = 8'b10011100;
DRAM[8829] = 8'b10101001;
DRAM[8830] = 8'b10110011;
DRAM[8831] = 8'b10111011;
DRAM[8832] = 8'b01100110;
DRAM[8833] = 8'b01101000;
DRAM[8834] = 8'b01100100;
DRAM[8835] = 8'b01011100;
DRAM[8836] = 8'b01010100;
DRAM[8837] = 8'b01001101;
DRAM[8838] = 8'b01010000;
DRAM[8839] = 8'b01111111;
DRAM[8840] = 8'b10011001;
DRAM[8841] = 8'b10101010;
DRAM[8842] = 8'b10110010;
DRAM[8843] = 8'b10110110;
DRAM[8844] = 8'b10110110;
DRAM[8845] = 8'b10110000;
DRAM[8846] = 8'b10011101;
DRAM[8847] = 8'b01111110;
DRAM[8848] = 8'b01010111;
DRAM[8849] = 8'b01011000;
DRAM[8850] = 8'b01100001;
DRAM[8851] = 8'b01100110;
DRAM[8852] = 8'b01101101;
DRAM[8853] = 8'b01101110;
DRAM[8854] = 8'b01100100;
DRAM[8855] = 8'b00111010;
DRAM[8856] = 8'b01111011;
DRAM[8857] = 8'b10011011;
DRAM[8858] = 8'b10001011;
DRAM[8859] = 8'b10000101;
DRAM[8860] = 8'b01101000;
DRAM[8861] = 8'b00110111;
DRAM[8862] = 8'b00110001;
DRAM[8863] = 8'b01101110;
DRAM[8864] = 8'b01011011;
DRAM[8865] = 8'b01001110;
DRAM[8866] = 8'b00111110;
DRAM[8867] = 8'b00101011;
DRAM[8868] = 8'b01011011;
DRAM[8869] = 8'b01001111;
DRAM[8870] = 8'b01000101;
DRAM[8871] = 8'b01100000;
DRAM[8872] = 8'b01101110;
DRAM[8873] = 8'b01110101;
DRAM[8874] = 8'b01101001;
DRAM[8875] = 8'b00101010;
DRAM[8876] = 8'b00101110;
DRAM[8877] = 8'b00101100;
DRAM[8878] = 8'b00101110;
DRAM[8879] = 8'b00101101;
DRAM[8880] = 8'b00110011;
DRAM[8881] = 8'b00100111;
DRAM[8882] = 8'b00100000;
DRAM[8883] = 8'b01101110;
DRAM[8884] = 8'b01101011;
DRAM[8885] = 8'b10101110;
DRAM[8886] = 8'b10101111;
DRAM[8887] = 8'b11000101;
DRAM[8888] = 8'b10111110;
DRAM[8889] = 8'b01101101;
DRAM[8890] = 8'b01110111;
DRAM[8891] = 8'b10001000;
DRAM[8892] = 8'b10001011;
DRAM[8893] = 8'b10010001;
DRAM[8894] = 8'b10010000;
DRAM[8895] = 8'b10001100;
DRAM[8896] = 8'b10000111;
DRAM[8897] = 8'b01111000;
DRAM[8898] = 8'b01110001;
DRAM[8899] = 8'b01111010;
DRAM[8900] = 8'b01111001;
DRAM[8901] = 8'b10100000;
DRAM[8902] = 8'b10100101;
DRAM[8903] = 8'b10001110;
DRAM[8904] = 8'b01111000;
DRAM[8905] = 8'b10000001;
DRAM[8906] = 8'b10000001;
DRAM[8907] = 8'b10000111;
DRAM[8908] = 8'b10100110;
DRAM[8909] = 8'b11010111;
DRAM[8910] = 8'b11001000;
DRAM[8911] = 8'b10100010;
DRAM[8912] = 8'b10001110;
DRAM[8913] = 8'b10000000;
DRAM[8914] = 8'b01110001;
DRAM[8915] = 8'b01011110;
DRAM[8916] = 8'b01001000;
DRAM[8917] = 8'b01001101;
DRAM[8918] = 8'b01001110;
DRAM[8919] = 8'b00111000;
DRAM[8920] = 8'b00101111;
DRAM[8921] = 8'b00110101;
DRAM[8922] = 8'b01000000;
DRAM[8923] = 8'b01101010;
DRAM[8924] = 8'b10100110;
DRAM[8925] = 8'b01010001;
DRAM[8926] = 8'b01010001;
DRAM[8927] = 8'b00110110;
DRAM[8928] = 8'b00110001;
DRAM[8929] = 8'b00110101;
DRAM[8930] = 8'b00110100;
DRAM[8931] = 8'b01000111;
DRAM[8932] = 8'b10000010;
DRAM[8933] = 8'b10000101;
DRAM[8934] = 8'b10010100;
DRAM[8935] = 8'b10011101;
DRAM[8936] = 8'b10011100;
DRAM[8937] = 8'b10011010;
DRAM[8938] = 8'b10011001;
DRAM[8939] = 8'b10010111;
DRAM[8940] = 8'b10010111;
DRAM[8941] = 8'b10011010;
DRAM[8942] = 8'b10011000;
DRAM[8943] = 8'b10011000;
DRAM[8944] = 8'b10010111;
DRAM[8945] = 8'b10011000;
DRAM[8946] = 8'b10010111;
DRAM[8947] = 8'b10010100;
DRAM[8948] = 8'b10010010;
DRAM[8949] = 8'b10001101;
DRAM[8950] = 8'b10001001;
DRAM[8951] = 8'b10001001;
DRAM[8952] = 8'b10000111;
DRAM[8953] = 8'b10001100;
DRAM[8954] = 8'b10011011;
DRAM[8955] = 8'b10101100;
DRAM[8956] = 8'b10110110;
DRAM[8957] = 8'b10111011;
DRAM[8958] = 8'b10111011;
DRAM[8959] = 8'b10111101;
DRAM[8960] = 8'b01100100;
DRAM[8961] = 8'b01100011;
DRAM[8962] = 8'b01100000;
DRAM[8963] = 8'b01011000;
DRAM[8964] = 8'b01010010;
DRAM[8965] = 8'b01001010;
DRAM[8966] = 8'b01001000;
DRAM[8967] = 8'b01111100;
DRAM[8968] = 8'b10011000;
DRAM[8969] = 8'b10101010;
DRAM[8970] = 8'b10110000;
DRAM[8971] = 8'b10110011;
DRAM[8972] = 8'b10110110;
DRAM[8973] = 8'b10110001;
DRAM[8974] = 8'b10011110;
DRAM[8975] = 8'b01111100;
DRAM[8976] = 8'b01010101;
DRAM[8977] = 8'b01010110;
DRAM[8978] = 8'b01011111;
DRAM[8979] = 8'b01101001;
DRAM[8980] = 8'b01101110;
DRAM[8981] = 8'b01101011;
DRAM[8982] = 8'b10000011;
DRAM[8983] = 8'b10010101;
DRAM[8984] = 8'b10011001;
DRAM[8985] = 8'b10000110;
DRAM[8986] = 8'b01001000;
DRAM[8987] = 8'b01001010;
DRAM[8988] = 8'b01001011;
DRAM[8989] = 8'b00101010;
DRAM[8990] = 8'b00110100;
DRAM[8991] = 8'b00110111;
DRAM[8992] = 8'b01111010;
DRAM[8993] = 8'b10000010;
DRAM[8994] = 8'b01101010;
DRAM[8995] = 8'b00110000;
DRAM[8996] = 8'b01000011;
DRAM[8997] = 8'b00111111;
DRAM[8998] = 8'b01101011;
DRAM[8999] = 8'b01011000;
DRAM[9000] = 8'b01101010;
DRAM[9001] = 8'b10000100;
DRAM[9002] = 8'b01010101;
DRAM[9003] = 8'b01000001;
DRAM[9004] = 8'b00101110;
DRAM[9005] = 8'b00110010;
DRAM[9006] = 8'b00101110;
DRAM[9007] = 8'b00110011;
DRAM[9008] = 8'b00101111;
DRAM[9009] = 8'b00100011;
DRAM[9010] = 8'b00111100;
DRAM[9011] = 8'b01111111;
DRAM[9012] = 8'b10011110;
DRAM[9013] = 8'b10101001;
DRAM[9014] = 8'b10111101;
DRAM[9015] = 8'b11001110;
DRAM[9016] = 8'b01100101;
DRAM[9017] = 8'b01101001;
DRAM[9018] = 8'b01111110;
DRAM[9019] = 8'b10001010;
DRAM[9020] = 8'b10010111;
DRAM[9021] = 8'b10010100;
DRAM[9022] = 8'b10010111;
DRAM[9023] = 8'b10010100;
DRAM[9024] = 8'b10010001;
DRAM[9025] = 8'b10010000;
DRAM[9026] = 8'b10001101;
DRAM[9027] = 8'b10010100;
DRAM[9028] = 8'b10011110;
DRAM[9029] = 8'b10100011;
DRAM[9030] = 8'b10011100;
DRAM[9031] = 8'b10010011;
DRAM[9032] = 8'b10000001;
DRAM[9033] = 8'b10000111;
DRAM[9034] = 8'b10000000;
DRAM[9035] = 8'b10000000;
DRAM[9036] = 8'b10100110;
DRAM[9037] = 8'b11010000;
DRAM[9038] = 8'b11010001;
DRAM[9039] = 8'b10101110;
DRAM[9040] = 8'b10011011;
DRAM[9041] = 8'b10001100;
DRAM[9042] = 8'b10000010;
DRAM[9043] = 8'b01111000;
DRAM[9044] = 8'b01100011;
DRAM[9045] = 8'b01101000;
DRAM[9046] = 8'b01011010;
DRAM[9047] = 8'b00111000;
DRAM[9048] = 8'b00101110;
DRAM[9049] = 8'b00110100;
DRAM[9050] = 8'b00111101;
DRAM[9051] = 8'b01101010;
DRAM[9052] = 8'b10101011;
DRAM[9053] = 8'b01011011;
DRAM[9054] = 8'b01001110;
DRAM[9055] = 8'b00110000;
DRAM[9056] = 8'b00110000;
DRAM[9057] = 8'b00111010;
DRAM[9058] = 8'b00101001;
DRAM[9059] = 8'b01010100;
DRAM[9060] = 8'b10001000;
DRAM[9061] = 8'b10000101;
DRAM[9062] = 8'b10011010;
DRAM[9063] = 8'b10011100;
DRAM[9064] = 8'b10011001;
DRAM[9065] = 8'b10011011;
DRAM[9066] = 8'b10010111;
DRAM[9067] = 8'b10010101;
DRAM[9068] = 8'b10011000;
DRAM[9069] = 8'b10011000;
DRAM[9070] = 8'b10010101;
DRAM[9071] = 8'b10010111;
DRAM[9072] = 8'b10010110;
DRAM[9073] = 8'b10010111;
DRAM[9074] = 8'b10010011;
DRAM[9075] = 8'b10010011;
DRAM[9076] = 8'b10001110;
DRAM[9077] = 8'b10001101;
DRAM[9078] = 8'b10001001;
DRAM[9079] = 8'b10000110;
DRAM[9080] = 8'b10010010;
DRAM[9081] = 8'b10101010;
DRAM[9082] = 8'b10111000;
DRAM[9083] = 8'b10111110;
DRAM[9084] = 8'b10111110;
DRAM[9085] = 8'b10111110;
DRAM[9086] = 8'b10111110;
DRAM[9087] = 8'b10111110;
DRAM[9088] = 8'b01100011;
DRAM[9089] = 8'b01011000;
DRAM[9090] = 8'b01010110;
DRAM[9091] = 8'b01010010;
DRAM[9092] = 8'b01001110;
DRAM[9093] = 8'b01000001;
DRAM[9094] = 8'b01000100;
DRAM[9095] = 8'b01111001;
DRAM[9096] = 8'b10010111;
DRAM[9097] = 8'b10101000;
DRAM[9098] = 8'b10110010;
DRAM[9099] = 8'b10110111;
DRAM[9100] = 8'b10110111;
DRAM[9101] = 8'b10110001;
DRAM[9102] = 8'b10011110;
DRAM[9103] = 8'b10000000;
DRAM[9104] = 8'b01010101;
DRAM[9105] = 8'b01010100;
DRAM[9106] = 8'b01011110;
DRAM[9107] = 8'b01100111;
DRAM[9108] = 8'b01101110;
DRAM[9109] = 8'b01101100;
DRAM[9110] = 8'b01110001;
DRAM[9111] = 8'b10000110;
DRAM[9112] = 8'b01110011;
DRAM[9113] = 8'b01011100;
DRAM[9114] = 8'b01011110;
DRAM[9115] = 8'b01010101;
DRAM[9116] = 8'b00110111;
DRAM[9117] = 8'b00101110;
DRAM[9118] = 8'b01001100;
DRAM[9119] = 8'b01100101;
DRAM[9120] = 8'b01011101;
DRAM[9121] = 8'b01001000;
DRAM[9122] = 8'b01001100;
DRAM[9123] = 8'b00101000;
DRAM[9124] = 8'b00111010;
DRAM[9125] = 8'b01001111;
DRAM[9126] = 8'b01000001;
DRAM[9127] = 8'b10001110;
DRAM[9128] = 8'b01001110;
DRAM[9129] = 8'b01100010;
DRAM[9130] = 8'b01011110;
DRAM[9131] = 8'b00101100;
DRAM[9132] = 8'b00101111;
DRAM[9133] = 8'b00101100;
DRAM[9134] = 8'b00101010;
DRAM[9135] = 8'b00110001;
DRAM[9136] = 8'b00110011;
DRAM[9137] = 8'b00100111;
DRAM[9138] = 8'b01110101;
DRAM[9139] = 8'b01101110;
DRAM[9140] = 8'b10110001;
DRAM[9141] = 8'b10111011;
DRAM[9142] = 8'b11001101;
DRAM[9143] = 8'b01010101;
DRAM[9144] = 8'b01100000;
DRAM[9145] = 8'b01110100;
DRAM[9146] = 8'b10000010;
DRAM[9147] = 8'b10001010;
DRAM[9148] = 8'b10010111;
DRAM[9149] = 8'b10011110;
DRAM[9150] = 8'b10100101;
DRAM[9151] = 8'b10100100;
DRAM[9152] = 8'b10100101;
DRAM[9153] = 8'b10100010;
DRAM[9154] = 8'b10100011;
DRAM[9155] = 8'b10101011;
DRAM[9156] = 8'b10101010;
DRAM[9157] = 8'b10100111;
DRAM[9158] = 8'b10100001;
DRAM[9159] = 8'b10010000;
DRAM[9160] = 8'b10001010;
DRAM[9161] = 8'b10001010;
DRAM[9162] = 8'b10000001;
DRAM[9163] = 8'b10000000;
DRAM[9164] = 8'b10011111;
DRAM[9165] = 8'b11001011;
DRAM[9166] = 8'b11010101;
DRAM[9167] = 8'b10111001;
DRAM[9168] = 8'b10100010;
DRAM[9169] = 8'b10011000;
DRAM[9170] = 8'b10001100;
DRAM[9171] = 8'b10000100;
DRAM[9172] = 8'b01111010;
DRAM[9173] = 8'b01110100;
DRAM[9174] = 8'b01100010;
DRAM[9175] = 8'b00111011;
DRAM[9176] = 8'b00101100;
DRAM[9177] = 8'b00110111;
DRAM[9178] = 8'b01000000;
DRAM[9179] = 8'b01100010;
DRAM[9180] = 8'b10101101;
DRAM[9181] = 8'b01100010;
DRAM[9182] = 8'b00111110;
DRAM[9183] = 8'b00111010;
DRAM[9184] = 8'b00101010;
DRAM[9185] = 8'b00110000;
DRAM[9186] = 8'b00101101;
DRAM[9187] = 8'b01101001;
DRAM[9188] = 8'b10001000;
DRAM[9189] = 8'b10001010;
DRAM[9190] = 8'b10011101;
DRAM[9191] = 8'b10011010;
DRAM[9192] = 8'b10011100;
DRAM[9193] = 8'b10010111;
DRAM[9194] = 8'b10010110;
DRAM[9195] = 8'b10010110;
DRAM[9196] = 8'b10011000;
DRAM[9197] = 8'b10010111;
DRAM[9198] = 8'b10010101;
DRAM[9199] = 8'b10010110;
DRAM[9200] = 8'b10010111;
DRAM[9201] = 8'b10010011;
DRAM[9202] = 8'b10010010;
DRAM[9203] = 8'b10010000;
DRAM[9204] = 8'b10001101;
DRAM[9205] = 8'b10001001;
DRAM[9206] = 8'b10000101;
DRAM[9207] = 8'b10010011;
DRAM[9208] = 8'b10110010;
DRAM[9209] = 8'b11000001;
DRAM[9210] = 8'b11000011;
DRAM[9211] = 8'b11000000;
DRAM[9212] = 8'b10111111;
DRAM[9213] = 8'b10111110;
DRAM[9214] = 8'b10111110;
DRAM[9215] = 8'b10111110;
DRAM[9216] = 8'b01011100;
DRAM[9217] = 8'b01011101;
DRAM[9218] = 8'b01010110;
DRAM[9219] = 8'b01010001;
DRAM[9220] = 8'b01001011;
DRAM[9221] = 8'b01000000;
DRAM[9222] = 8'b01000100;
DRAM[9223] = 8'b01111000;
DRAM[9224] = 8'b10010101;
DRAM[9225] = 8'b10101001;
DRAM[9226] = 8'b10110010;
DRAM[9227] = 8'b10110100;
DRAM[9228] = 8'b10110110;
DRAM[9229] = 8'b10110001;
DRAM[9230] = 8'b10011101;
DRAM[9231] = 8'b01111110;
DRAM[9232] = 8'b01010110;
DRAM[9233] = 8'b01010011;
DRAM[9234] = 8'b01011100;
DRAM[9235] = 8'b01100101;
DRAM[9236] = 8'b01101110;
DRAM[9237] = 8'b01111100;
DRAM[9238] = 8'b10001011;
DRAM[9239] = 8'b10001000;
DRAM[9240] = 8'b10011101;
DRAM[9241] = 8'b01110010;
DRAM[9242] = 8'b01101110;
DRAM[9243] = 8'b00111101;
DRAM[9244] = 8'b00111111;
DRAM[9245] = 8'b01001000;
DRAM[9246] = 8'b01010110;
DRAM[9247] = 8'b01110000;
DRAM[9248] = 8'b01100000;
DRAM[9249] = 8'b01100110;
DRAM[9250] = 8'b00101101;
DRAM[9251] = 8'b00101000;
DRAM[9252] = 8'b00110001;
DRAM[9253] = 8'b01011010;
DRAM[9254] = 8'b01100010;
DRAM[9255] = 8'b01100100;
DRAM[9256] = 8'b01111001;
DRAM[9257] = 8'b10000100;
DRAM[9258] = 8'b01010100;
DRAM[9259] = 8'b01010001;
DRAM[9260] = 8'b00110110;
DRAM[9261] = 8'b00110001;
DRAM[9262] = 8'b00101100;
DRAM[9263] = 8'b00110001;
DRAM[9264] = 8'b00101101;
DRAM[9265] = 8'b01010000;
DRAM[9266] = 8'b01111010;
DRAM[9267] = 8'b10011010;
DRAM[9268] = 8'b10111000;
DRAM[9269] = 8'b11000100;
DRAM[9270] = 8'b01111001;
DRAM[9271] = 8'b01000101;
DRAM[9272] = 8'b01101000;
DRAM[9273] = 8'b01111000;
DRAM[9274] = 8'b10000011;
DRAM[9275] = 8'b10001010;
DRAM[9276] = 8'b10010110;
DRAM[9277] = 8'b10011110;
DRAM[9278] = 8'b10100101;
DRAM[9279] = 8'b10101000;
DRAM[9280] = 8'b10101100;
DRAM[9281] = 8'b10101110;
DRAM[9282] = 8'b10101110;
DRAM[9283] = 8'b10101001;
DRAM[9284] = 8'b10101011;
DRAM[9285] = 8'b10101011;
DRAM[9286] = 8'b10011110;
DRAM[9287] = 8'b10010010;
DRAM[9288] = 8'b10010001;
DRAM[9289] = 8'b10000111;
DRAM[9290] = 8'b10000010;
DRAM[9291] = 8'b10000001;
DRAM[9292] = 8'b10010110;
DRAM[9293] = 8'b11001011;
DRAM[9294] = 8'b11011001;
DRAM[9295] = 8'b10110110;
DRAM[9296] = 8'b10101100;
DRAM[9297] = 8'b10011001;
DRAM[9298] = 8'b10001101;
DRAM[9299] = 8'b10000111;
DRAM[9300] = 8'b10000010;
DRAM[9301] = 8'b01110111;
DRAM[9302] = 8'b01100110;
DRAM[9303] = 8'b00111011;
DRAM[9304] = 8'b00110001;
DRAM[9305] = 8'b00111111;
DRAM[9306] = 8'b01000001;
DRAM[9307] = 8'b01010100;
DRAM[9308] = 8'b10101010;
DRAM[9309] = 8'b01100110;
DRAM[9310] = 8'b00110101;
DRAM[9311] = 8'b00110011;
DRAM[9312] = 8'b00101110;
DRAM[9313] = 8'b00110010;
DRAM[9314] = 8'b00110111;
DRAM[9315] = 8'b01111111;
DRAM[9316] = 8'b10000110;
DRAM[9317] = 8'b10010001;
DRAM[9318] = 8'b10011111;
DRAM[9319] = 8'b10011001;
DRAM[9320] = 8'b10011010;
DRAM[9321] = 8'b10011000;
DRAM[9322] = 8'b10010110;
DRAM[9323] = 8'b10010110;
DRAM[9324] = 8'b10011000;
DRAM[9325] = 8'b10010111;
DRAM[9326] = 8'b10010101;
DRAM[9327] = 8'b10010101;
DRAM[9328] = 8'b10010010;
DRAM[9329] = 8'b10010001;
DRAM[9330] = 8'b10010000;
DRAM[9331] = 8'b10001011;
DRAM[9332] = 8'b10001010;
DRAM[9333] = 8'b10000110;
DRAM[9334] = 8'b10001111;
DRAM[9335] = 8'b10110010;
DRAM[9336] = 8'b11000001;
DRAM[9337] = 8'b11000110;
DRAM[9338] = 8'b11000100;
DRAM[9339] = 8'b11000001;
DRAM[9340] = 8'b10111110;
DRAM[9341] = 8'b10111101;
DRAM[9342] = 8'b10111111;
DRAM[9343] = 8'b11000001;
DRAM[9344] = 8'b01010110;
DRAM[9345] = 8'b01010110;
DRAM[9346] = 8'b01010001;
DRAM[9347] = 8'b01001111;
DRAM[9348] = 8'b01001000;
DRAM[9349] = 8'b00111111;
DRAM[9350] = 8'b01000010;
DRAM[9351] = 8'b01111000;
DRAM[9352] = 8'b10010111;
DRAM[9353] = 8'b10100111;
DRAM[9354] = 8'b10110000;
DRAM[9355] = 8'b10110011;
DRAM[9356] = 8'b10110110;
DRAM[9357] = 8'b10110000;
DRAM[9358] = 8'b10011100;
DRAM[9359] = 8'b01111110;
DRAM[9360] = 8'b01010010;
DRAM[9361] = 8'b01010010;
DRAM[9362] = 8'b01011100;
DRAM[9363] = 8'b01101110;
DRAM[9364] = 8'b10000001;
DRAM[9365] = 8'b10000010;
DRAM[9366] = 8'b10000000;
DRAM[9367] = 8'b01111010;
DRAM[9368] = 8'b01001110;
DRAM[9369] = 8'b01001000;
DRAM[9370] = 8'b01000100;
DRAM[9371] = 8'b00111101;
DRAM[9372] = 8'b01000011;
DRAM[9373] = 8'b01010100;
DRAM[9374] = 8'b01100100;
DRAM[9375] = 8'b01110000;
DRAM[9376] = 8'b01111111;
DRAM[9377] = 8'b00110101;
DRAM[9378] = 8'b00110010;
DRAM[9379] = 8'b00101100;
DRAM[9380] = 8'b00101111;
DRAM[9381] = 8'b00110011;
DRAM[9382] = 8'b01001010;
DRAM[9383] = 8'b01100011;
DRAM[9384] = 8'b01000011;
DRAM[9385] = 8'b00100111;
DRAM[9386] = 8'b01111010;
DRAM[9387] = 8'b01101110;
DRAM[9388] = 8'b00111011;
DRAM[9389] = 8'b00101011;
DRAM[9390] = 8'b00101111;
DRAM[9391] = 8'b00101011;
DRAM[9392] = 8'b00101011;
DRAM[9393] = 8'b10000001;
DRAM[9394] = 8'b01110100;
DRAM[9395] = 8'b10111010;
DRAM[9396] = 8'b11000011;
DRAM[9397] = 8'b10101000;
DRAM[9398] = 8'b00101000;
DRAM[9399] = 8'b01001110;
DRAM[9400] = 8'b01110010;
DRAM[9401] = 8'b01111010;
DRAM[9402] = 8'b10000000;
DRAM[9403] = 8'b10001011;
DRAM[9404] = 8'b10010101;
DRAM[9405] = 8'b10011011;
DRAM[9406] = 8'b10100101;
DRAM[9407] = 8'b10101100;
DRAM[9408] = 8'b10110001;
DRAM[9409] = 8'b10101111;
DRAM[9410] = 8'b10110000;
DRAM[9411] = 8'b10110000;
DRAM[9412] = 8'b10110000;
DRAM[9413] = 8'b10101010;
DRAM[9414] = 8'b10100000;
DRAM[9415] = 8'b10010101;
DRAM[9416] = 8'b10010001;
DRAM[9417] = 8'b10001001;
DRAM[9418] = 8'b10000011;
DRAM[9419] = 8'b10000001;
DRAM[9420] = 8'b10010100;
DRAM[9421] = 8'b11000110;
DRAM[9422] = 8'b11011010;
DRAM[9423] = 8'b10111011;
DRAM[9424] = 8'b10100101;
DRAM[9425] = 8'b10011110;
DRAM[9426] = 8'b10010000;
DRAM[9427] = 8'b10000111;
DRAM[9428] = 8'b10000000;
DRAM[9429] = 8'b01111101;
DRAM[9430] = 8'b01100101;
DRAM[9431] = 8'b00111001;
DRAM[9432] = 8'b00110101;
DRAM[9433] = 8'b01000010;
DRAM[9434] = 8'b01000000;
DRAM[9435] = 8'b01000010;
DRAM[9436] = 8'b10100101;
DRAM[9437] = 8'b10001010;
DRAM[9438] = 8'b00101111;
DRAM[9439] = 8'b00101011;
DRAM[9440] = 8'b00110011;
DRAM[9441] = 8'b00101010;
DRAM[9442] = 8'b01000110;
DRAM[9443] = 8'b10000111;
DRAM[9444] = 8'b10000111;
DRAM[9445] = 8'b10011011;
DRAM[9446] = 8'b10011110;
DRAM[9447] = 8'b10011010;
DRAM[9448] = 8'b10011010;
DRAM[9449] = 8'b10011000;
DRAM[9450] = 8'b10010111;
DRAM[9451] = 8'b10011010;
DRAM[9452] = 8'b10010100;
DRAM[9453] = 8'b10010101;
DRAM[9454] = 8'b10010010;
DRAM[9455] = 8'b10010010;
DRAM[9456] = 8'b10010010;
DRAM[9457] = 8'b10001111;
DRAM[9458] = 8'b10001110;
DRAM[9459] = 8'b10001011;
DRAM[9460] = 8'b10000101;
DRAM[9461] = 8'b10001001;
DRAM[9462] = 8'b10101110;
DRAM[9463] = 8'b10111111;
DRAM[9464] = 8'b11000010;
DRAM[9465] = 8'b11000100;
DRAM[9466] = 8'b11000010;
DRAM[9467] = 8'b11000010;
DRAM[9468] = 8'b10111111;
DRAM[9469] = 8'b11000000;
DRAM[9470] = 8'b11000100;
DRAM[9471] = 8'b11000110;
DRAM[9472] = 8'b01010000;
DRAM[9473] = 8'b01001101;
DRAM[9474] = 8'b01001110;
DRAM[9475] = 8'b01001010;
DRAM[9476] = 8'b01001000;
DRAM[9477] = 8'b00111101;
DRAM[9478] = 8'b00111101;
DRAM[9479] = 8'b01110111;
DRAM[9480] = 8'b10010110;
DRAM[9481] = 8'b10101000;
DRAM[9482] = 8'b10110010;
DRAM[9483] = 8'b10110011;
DRAM[9484] = 8'b10110011;
DRAM[9485] = 8'b10101111;
DRAM[9486] = 8'b10011011;
DRAM[9487] = 8'b01111010;
DRAM[9488] = 8'b01010101;
DRAM[9489] = 8'b01010101;
DRAM[9490] = 8'b01011101;
DRAM[9491] = 8'b01100110;
DRAM[9492] = 8'b01101111;
DRAM[9493] = 8'b01110100;
DRAM[9494] = 8'b01101011;
DRAM[9495] = 8'b01010110;
DRAM[9496] = 8'b01011011;
DRAM[9497] = 8'b01011101;
DRAM[9498] = 8'b01001010;
DRAM[9499] = 8'b01000010;
DRAM[9500] = 8'b01100110;
DRAM[9501] = 8'b01000000;
DRAM[9502] = 8'b01110110;
DRAM[9503] = 8'b01101110;
DRAM[9504] = 8'b01001000;
DRAM[9505] = 8'b00110010;
DRAM[9506] = 8'b00101111;
DRAM[9507] = 8'b00110010;
DRAM[9508] = 8'b00101111;
DRAM[9509] = 8'b00110001;
DRAM[9510] = 8'b00110001;
DRAM[9511] = 8'b00111101;
DRAM[9512] = 8'b00111100;
DRAM[9513] = 8'b00100101;
DRAM[9514] = 8'b01111010;
DRAM[9515] = 8'b10000101;
DRAM[9516] = 8'b00111111;
DRAM[9517] = 8'b00101001;
DRAM[9518] = 8'b00101000;
DRAM[9519] = 8'b00100110;
DRAM[9520] = 8'b01001100;
DRAM[9521] = 8'b01111101;
DRAM[9522] = 8'b10011110;
DRAM[9523] = 8'b10111011;
DRAM[9524] = 8'b11000110;
DRAM[9525] = 8'b00110011;
DRAM[9526] = 8'b00110010;
DRAM[9527] = 8'b01010110;
DRAM[9528] = 8'b01110101;
DRAM[9529] = 8'b01111101;
DRAM[9530] = 8'b10000001;
DRAM[9531] = 8'b10000111;
DRAM[9532] = 8'b10010001;
DRAM[9533] = 8'b10010110;
DRAM[9534] = 8'b10011110;
DRAM[9535] = 8'b10101100;
DRAM[9536] = 8'b10110000;
DRAM[9537] = 8'b10110010;
DRAM[9538] = 8'b10110100;
DRAM[9539] = 8'b10101110;
DRAM[9540] = 8'b10101101;
DRAM[9541] = 8'b10101000;
DRAM[9542] = 8'b10011101;
DRAM[9543] = 8'b10010011;
DRAM[9544] = 8'b10010010;
DRAM[9545] = 8'b10001100;
DRAM[9546] = 8'b10000010;
DRAM[9547] = 8'b10000011;
DRAM[9548] = 8'b10010000;
DRAM[9549] = 8'b11000000;
DRAM[9550] = 8'b11011101;
DRAM[9551] = 8'b10111101;
DRAM[9552] = 8'b10100100;
DRAM[9553] = 8'b10011110;
DRAM[9554] = 8'b10010011;
DRAM[9555] = 8'b10001001;
DRAM[9556] = 8'b10000011;
DRAM[9557] = 8'b01111110;
DRAM[9558] = 8'b01011011;
DRAM[9559] = 8'b00110111;
DRAM[9560] = 8'b00110011;
DRAM[9561] = 8'b00111101;
DRAM[9562] = 8'b00111100;
DRAM[9563] = 8'b00110100;
DRAM[9564] = 8'b10100111;
DRAM[9565] = 8'b10011011;
DRAM[9566] = 8'b00100010;
DRAM[9567] = 8'b00110001;
DRAM[9568] = 8'b00110111;
DRAM[9569] = 8'b00101100;
DRAM[9570] = 8'b01011010;
DRAM[9571] = 8'b10001011;
DRAM[9572] = 8'b10001100;
DRAM[9573] = 8'b10100001;
DRAM[9574] = 8'b10011101;
DRAM[9575] = 8'b10010111;
DRAM[9576] = 8'b10011010;
DRAM[9577] = 8'b10011010;
DRAM[9578] = 8'b10010110;
DRAM[9579] = 8'b10010110;
DRAM[9580] = 8'b10010110;
DRAM[9581] = 8'b10010010;
DRAM[9582] = 8'b10010011;
DRAM[9583] = 8'b10010010;
DRAM[9584] = 8'b10010010;
DRAM[9585] = 8'b10010001;
DRAM[9586] = 8'b10001100;
DRAM[9587] = 8'b10000111;
DRAM[9588] = 8'b10000001;
DRAM[9589] = 8'b10100011;
DRAM[9590] = 8'b10111101;
DRAM[9591] = 8'b11000011;
DRAM[9592] = 8'b11000001;
DRAM[9593] = 8'b11000010;
DRAM[9594] = 8'b11000010;
DRAM[9595] = 8'b11000010;
DRAM[9596] = 8'b11000010;
DRAM[9597] = 8'b11000111;
DRAM[9598] = 8'b11001100;
DRAM[9599] = 8'b11001100;
DRAM[9600] = 8'b01001110;
DRAM[9601] = 8'b01001010;
DRAM[9602] = 8'b01001010;
DRAM[9603] = 8'b01000110;
DRAM[9604] = 8'b01000100;
DRAM[9605] = 8'b00111001;
DRAM[9606] = 8'b00111111;
DRAM[9607] = 8'b01110101;
DRAM[9608] = 8'b10010111;
DRAM[9609] = 8'b10101000;
DRAM[9610] = 8'b10101101;
DRAM[9611] = 8'b10101110;
DRAM[9612] = 8'b10110001;
DRAM[9613] = 8'b10101100;
DRAM[9614] = 8'b10011011;
DRAM[9615] = 8'b01111111;
DRAM[9616] = 8'b01010101;
DRAM[9617] = 8'b01010010;
DRAM[9618] = 8'b01100100;
DRAM[9619] = 8'b01100011;
DRAM[9620] = 8'b01101011;
DRAM[9621] = 8'b01101111;
DRAM[9622] = 8'b01100111;
DRAM[9623] = 8'b10000111;
DRAM[9624] = 8'b01010110;
DRAM[9625] = 8'b01100000;
DRAM[9626] = 8'b01001111;
DRAM[9627] = 8'b01100100;
DRAM[9628] = 8'b00111100;
DRAM[9629] = 8'b00110111;
DRAM[9630] = 8'b01010001;
DRAM[9631] = 8'b01100011;
DRAM[9632] = 8'b00111110;
DRAM[9633] = 8'b00111100;
DRAM[9634] = 8'b00110100;
DRAM[9635] = 8'b00110001;
DRAM[9636] = 8'b00110001;
DRAM[9637] = 8'b00101111;
DRAM[9638] = 8'b00110110;
DRAM[9639] = 8'b00111111;
DRAM[9640] = 8'b00110101;
DRAM[9641] = 8'b00101111;
DRAM[9642] = 8'b01110100;
DRAM[9643] = 8'b01110101;
DRAM[9644] = 8'b10000100;
DRAM[9645] = 8'b00101110;
DRAM[9646] = 8'b00100100;
DRAM[9647] = 8'b00100110;
DRAM[9648] = 8'b01111011;
DRAM[9649] = 8'b01110011;
DRAM[9650] = 8'b11000011;
DRAM[9651] = 8'b11001011;
DRAM[9652] = 8'b01100010;
DRAM[9653] = 8'b00110001;
DRAM[9654] = 8'b00110100;
DRAM[9655] = 8'b01010100;
DRAM[9656] = 8'b01110100;
DRAM[9657] = 8'b01111010;
DRAM[9658] = 8'b10000010;
DRAM[9659] = 8'b10001001;
DRAM[9660] = 8'b10010000;
DRAM[9661] = 8'b10010111;
DRAM[9662] = 8'b10011011;
DRAM[9663] = 8'b10100001;
DRAM[9664] = 8'b10100111;
DRAM[9665] = 8'b10110000;
DRAM[9666] = 8'b10110010;
DRAM[9667] = 8'b10101100;
DRAM[9668] = 8'b10101010;
DRAM[9669] = 8'b10100001;
DRAM[9670] = 8'b10011001;
DRAM[9671] = 8'b10001110;
DRAM[9672] = 8'b10001100;
DRAM[9673] = 8'b10001000;
DRAM[9674] = 8'b01111100;
DRAM[9675] = 8'b10000000;
DRAM[9676] = 8'b10010000;
DRAM[9677] = 8'b10110000;
DRAM[9678] = 8'b11011100;
DRAM[9679] = 8'b10111110;
DRAM[9680] = 8'b10100011;
DRAM[9681] = 8'b10011100;
DRAM[9682] = 8'b10010111;
DRAM[9683] = 8'b10001100;
DRAM[9684] = 8'b10000011;
DRAM[9685] = 8'b01111100;
DRAM[9686] = 8'b01010001;
DRAM[9687] = 8'b00101111;
DRAM[9688] = 8'b00110111;
DRAM[9689] = 8'b00111111;
DRAM[9690] = 8'b00111000;
DRAM[9691] = 8'b00101110;
DRAM[9692] = 8'b10101110;
DRAM[9693] = 8'b10010010;
DRAM[9694] = 8'b00111001;
DRAM[9695] = 8'b00101010;
DRAM[9696] = 8'b00110111;
DRAM[9697] = 8'b00110100;
DRAM[9698] = 8'b01110010;
DRAM[9699] = 8'b10001001;
DRAM[9700] = 8'b10011001;
DRAM[9701] = 8'b10101011;
DRAM[9702] = 8'b10011100;
DRAM[9703] = 8'b10011011;
DRAM[9704] = 8'b10011011;
DRAM[9705] = 8'b10011000;
DRAM[9706] = 8'b10010110;
DRAM[9707] = 8'b10010100;
DRAM[9708] = 8'b10010001;
DRAM[9709] = 8'b10010010;
DRAM[9710] = 8'b10010000;
DRAM[9711] = 8'b10010000;
DRAM[9712] = 8'b10001111;
DRAM[9713] = 8'b10001110;
DRAM[9714] = 8'b10001010;
DRAM[9715] = 8'b10000011;
DRAM[9716] = 8'b10010000;
DRAM[9717] = 8'b10111001;
DRAM[9718] = 8'b11000011;
DRAM[9719] = 8'b11000010;
DRAM[9720] = 8'b11000000;
DRAM[9721] = 8'b11000001;
DRAM[9722] = 8'b11000010;
DRAM[9723] = 8'b11000111;
DRAM[9724] = 8'b11001010;
DRAM[9725] = 8'b11001101;
DRAM[9726] = 8'b11001100;
DRAM[9727] = 8'b11001011;
DRAM[9728] = 8'b01001011;
DRAM[9729] = 8'b01001011;
DRAM[9730] = 8'b01001100;
DRAM[9731] = 8'b01000110;
DRAM[9732] = 8'b01000100;
DRAM[9733] = 8'b00110111;
DRAM[9734] = 8'b00111110;
DRAM[9735] = 8'b01110101;
DRAM[9736] = 8'b10010101;
DRAM[9737] = 8'b10100101;
DRAM[9738] = 8'b10101110;
DRAM[9739] = 8'b10101101;
DRAM[9740] = 8'b10110011;
DRAM[9741] = 8'b10101100;
DRAM[9742] = 8'b10011010;
DRAM[9743] = 8'b01111110;
DRAM[9744] = 8'b01001111;
DRAM[9745] = 8'b01001110;
DRAM[9746] = 8'b01111111;
DRAM[9747] = 8'b01100000;
DRAM[9748] = 8'b10000001;
DRAM[9749] = 8'b10001101;
DRAM[9750] = 8'b01101011;
DRAM[9751] = 8'b00110000;
DRAM[9752] = 8'b01101110;
DRAM[9753] = 8'b01110110;
DRAM[9754] = 8'b01101100;
DRAM[9755] = 8'b00110000;
DRAM[9756] = 8'b01010110;
DRAM[9757] = 8'b01000100;
DRAM[9758] = 8'b01100100;
DRAM[9759] = 8'b01101110;
DRAM[9760] = 8'b01100110;
DRAM[9761] = 8'b00110101;
DRAM[9762] = 8'b00111010;
DRAM[9763] = 8'b00110110;
DRAM[9764] = 8'b00101000;
DRAM[9765] = 8'b00101110;
DRAM[9766] = 8'b00111010;
DRAM[9767] = 8'b01001101;
DRAM[9768] = 8'b00111011;
DRAM[9769] = 8'b01001110;
DRAM[9770] = 8'b10001001;
DRAM[9771] = 8'b01100100;
DRAM[9772] = 8'b01110110;
DRAM[9773] = 8'b01010100;
DRAM[9774] = 8'b00100000;
DRAM[9775] = 8'b01000010;
DRAM[9776] = 8'b01111100;
DRAM[9777] = 8'b10010101;
DRAM[9778] = 8'b11001010;
DRAM[9779] = 8'b10101001;
DRAM[9780] = 8'b00100001;
DRAM[9781] = 8'b00110010;
DRAM[9782] = 8'b00111000;
DRAM[9783] = 8'b01010010;
DRAM[9784] = 8'b01101010;
DRAM[9785] = 8'b01111000;
DRAM[9786] = 8'b10000011;
DRAM[9787] = 8'b10000100;
DRAM[9788] = 8'b10001101;
DRAM[9789] = 8'b10010100;
DRAM[9790] = 8'b10011011;
DRAM[9791] = 8'b10100000;
DRAM[9792] = 8'b10100100;
DRAM[9793] = 8'b10101101;
DRAM[9794] = 8'b10101010;
DRAM[9795] = 8'b10101010;
DRAM[9796] = 8'b10101001;
DRAM[9797] = 8'b10100001;
DRAM[9798] = 8'b10010111;
DRAM[9799] = 8'b10000110;
DRAM[9800] = 8'b10000101;
DRAM[9801] = 8'b10000011;
DRAM[9802] = 8'b01111101;
DRAM[9803] = 8'b01111110;
DRAM[9804] = 8'b10001001;
DRAM[9805] = 8'b10101111;
DRAM[9806] = 8'b11010111;
DRAM[9807] = 8'b11000110;
DRAM[9808] = 8'b10100001;
DRAM[9809] = 8'b10011011;
DRAM[9810] = 8'b10010010;
DRAM[9811] = 8'b10001011;
DRAM[9812] = 8'b10000001;
DRAM[9813] = 8'b01111001;
DRAM[9814] = 8'b01000101;
DRAM[9815] = 8'b00101110;
DRAM[9816] = 8'b00111100;
DRAM[9817] = 8'b01000010;
DRAM[9818] = 8'b00111111;
DRAM[9819] = 8'b00101001;
DRAM[9820] = 8'b10100000;
DRAM[9821] = 8'b10001000;
DRAM[9822] = 8'b01010001;
DRAM[9823] = 8'b00101101;
DRAM[9824] = 8'b00110011;
DRAM[9825] = 8'b00111001;
DRAM[9826] = 8'b10000110;
DRAM[9827] = 8'b10001000;
DRAM[9828] = 8'b10011110;
DRAM[9829] = 8'b10011111;
DRAM[9830] = 8'b10011100;
DRAM[9831] = 8'b10011100;
DRAM[9832] = 8'b10011011;
DRAM[9833] = 8'b10010101;
DRAM[9834] = 8'b10010110;
DRAM[9835] = 8'b10010100;
DRAM[9836] = 8'b10010010;
DRAM[9837] = 8'b10010011;
DRAM[9838] = 8'b10010010;
DRAM[9839] = 8'b10001111;
DRAM[9840] = 8'b10001011;
DRAM[9841] = 8'b10001110;
DRAM[9842] = 8'b10001001;
DRAM[9843] = 8'b10000100;
DRAM[9844] = 8'b10101010;
DRAM[9845] = 8'b11000000;
DRAM[9846] = 8'b11000010;
DRAM[9847] = 8'b11000001;
DRAM[9848] = 8'b11000001;
DRAM[9849] = 8'b11000010;
DRAM[9850] = 8'b11000111;
DRAM[9851] = 8'b11001101;
DRAM[9852] = 8'b11010010;
DRAM[9853] = 8'b11001111;
DRAM[9854] = 8'b11001011;
DRAM[9855] = 8'b11001010;
DRAM[9856] = 8'b01001110;
DRAM[9857] = 8'b01001101;
DRAM[9858] = 8'b01001110;
DRAM[9859] = 8'b01000101;
DRAM[9860] = 8'b00111110;
DRAM[9861] = 8'b00110110;
DRAM[9862] = 8'b00111000;
DRAM[9863] = 8'b01110010;
DRAM[9864] = 8'b10010101;
DRAM[9865] = 8'b10101000;
DRAM[9866] = 8'b10101101;
DRAM[9867] = 8'b10101100;
DRAM[9868] = 8'b10110000;
DRAM[9869] = 8'b10101100;
DRAM[9870] = 8'b10011100;
DRAM[9871] = 8'b01111111;
DRAM[9872] = 8'b01010000;
DRAM[9873] = 8'b01001101;
DRAM[9874] = 8'b01101110;
DRAM[9875] = 8'b10000011;
DRAM[9876] = 8'b01111011;
DRAM[9877] = 8'b01111000;
DRAM[9878] = 8'b01011000;
DRAM[9879] = 8'b01011010;
DRAM[9880] = 8'b01101110;
DRAM[9881] = 8'b01100000;
DRAM[9882] = 8'b01000110;
DRAM[9883] = 8'b01000101;
DRAM[9884] = 8'b01100000;
DRAM[9885] = 8'b01011010;
DRAM[9886] = 8'b01111111;
DRAM[9887] = 8'b10000010;
DRAM[9888] = 8'b01100111;
DRAM[9889] = 8'b00101110;
DRAM[9890] = 8'b00111001;
DRAM[9891] = 8'b00110001;
DRAM[9892] = 8'b00100111;
DRAM[9893] = 8'b00101110;
DRAM[9894] = 8'b01001110;
DRAM[9895] = 8'b01100011;
DRAM[9896] = 8'b01000111;
DRAM[9897] = 8'b01101111;
DRAM[9898] = 8'b10010010;
DRAM[9899] = 8'b10010110;
DRAM[9900] = 8'b00111011;
DRAM[9901] = 8'b00111110;
DRAM[9902] = 8'b00011110;
DRAM[9903] = 8'b01110010;
DRAM[9904] = 8'b01110010;
DRAM[9905] = 8'b10111000;
DRAM[9906] = 8'b11001001;
DRAM[9907] = 8'b00101110;
DRAM[9908] = 8'b00100011;
DRAM[9909] = 8'b00111010;
DRAM[9910] = 8'b01000100;
DRAM[9911] = 8'b01001111;
DRAM[9912] = 8'b01101100;
DRAM[9913] = 8'b01111100;
DRAM[9914] = 8'b01111111;
DRAM[9915] = 8'b10000101;
DRAM[9916] = 8'b10001010;
DRAM[9917] = 8'b10010010;
DRAM[9918] = 8'b10011000;
DRAM[9919] = 8'b10011010;
DRAM[9920] = 8'b10100000;
DRAM[9921] = 8'b10100011;
DRAM[9922] = 8'b10100111;
DRAM[9923] = 8'b10100111;
DRAM[9924] = 8'b10100011;
DRAM[9925] = 8'b10100010;
DRAM[9926] = 8'b10010010;
DRAM[9927] = 8'b10000110;
DRAM[9928] = 8'b10000010;
DRAM[9929] = 8'b01111111;
DRAM[9930] = 8'b01111100;
DRAM[9931] = 8'b01111011;
DRAM[9932] = 8'b10000111;
DRAM[9933] = 8'b10100111;
DRAM[9934] = 8'b11010011;
DRAM[9935] = 8'b11011011;
DRAM[9936] = 8'b10011010;
DRAM[9937] = 8'b10011001;
DRAM[9938] = 8'b10010001;
DRAM[9939] = 8'b10001000;
DRAM[9940] = 8'b10000001;
DRAM[9941] = 8'b01101110;
DRAM[9942] = 8'b00111001;
DRAM[9943] = 8'b00110000;
DRAM[9944] = 8'b00110111;
DRAM[9945] = 8'b01000010;
DRAM[9946] = 8'b01000000;
DRAM[9947] = 8'b00101000;
DRAM[9948] = 8'b10010010;
DRAM[9949] = 8'b10011110;
DRAM[9950] = 8'b01010100;
DRAM[9951] = 8'b00101100;
DRAM[9952] = 8'b00101011;
DRAM[9953] = 8'b01010010;
DRAM[9954] = 8'b10001100;
DRAM[9955] = 8'b10001001;
DRAM[9956] = 8'b10011110;
DRAM[9957] = 8'b10011111;
DRAM[9958] = 8'b10011011;
DRAM[9959] = 8'b10010111;
DRAM[9960] = 8'b10011010;
DRAM[9961] = 8'b10010111;
DRAM[9962] = 8'b10010101;
DRAM[9963] = 8'b10010101;
DRAM[9964] = 8'b10010011;
DRAM[9965] = 8'b10010011;
DRAM[9966] = 8'b10010001;
DRAM[9967] = 8'b10010010;
DRAM[9968] = 8'b10001100;
DRAM[9969] = 8'b10001011;
DRAM[9970] = 8'b10000110;
DRAM[9971] = 8'b10010110;
DRAM[9972] = 8'b10111010;
DRAM[9973] = 8'b11000100;
DRAM[9974] = 8'b11000001;
DRAM[9975] = 8'b11000001;
DRAM[9976] = 8'b11000010;
DRAM[9977] = 8'b11000111;
DRAM[9978] = 8'b11001111;
DRAM[9979] = 8'b11010000;
DRAM[9980] = 8'b11010001;
DRAM[9981] = 8'b11010000;
DRAM[9982] = 8'b11001101;
DRAM[9983] = 8'b11001101;
DRAM[9984] = 8'b01001110;
DRAM[9985] = 8'b01001110;
DRAM[9986] = 8'b01001100;
DRAM[9987] = 8'b01001000;
DRAM[9988] = 8'b00111100;
DRAM[9989] = 8'b00110011;
DRAM[9990] = 8'b00110100;
DRAM[9991] = 8'b01110010;
DRAM[9992] = 8'b10010101;
DRAM[9993] = 8'b10100110;
DRAM[9994] = 8'b10101101;
DRAM[9995] = 8'b10110000;
DRAM[9996] = 8'b10110011;
DRAM[9997] = 8'b10101101;
DRAM[9998] = 8'b10011100;
DRAM[9999] = 8'b01111111;
DRAM[10000] = 8'b01010000;
DRAM[10001] = 8'b01001101;
DRAM[10002] = 8'b01011000;
DRAM[10003] = 8'b01110000;
DRAM[10004] = 8'b01110110;
DRAM[10005] = 8'b10000000;
DRAM[10006] = 8'b01011100;
DRAM[10007] = 8'b01011000;
DRAM[10008] = 8'b01010101;
DRAM[10009] = 8'b01100100;
DRAM[10010] = 8'b01001111;
DRAM[10011] = 8'b01010100;
DRAM[10012] = 8'b01101001;
DRAM[10013] = 8'b01000011;
DRAM[10014] = 8'b01011111;
DRAM[10015] = 8'b10010101;
DRAM[10016] = 8'b01001010;
DRAM[10017] = 8'b00101011;
DRAM[10018] = 8'b00101110;
DRAM[10019] = 8'b00111001;
DRAM[10020] = 8'b00110001;
DRAM[10021] = 8'b00101111;
DRAM[10022] = 8'b01001101;
DRAM[10023] = 8'b01001110;
DRAM[10024] = 8'b10000000;
DRAM[10025] = 8'b01100000;
DRAM[10026] = 8'b01001010;
DRAM[10027] = 8'b01000000;
DRAM[10028] = 8'b00101001;
DRAM[10029] = 8'b00101000;
DRAM[10030] = 8'b00111101;
DRAM[10031] = 8'b01111110;
DRAM[10032] = 8'b10001110;
DRAM[10033] = 8'b10110111;
DRAM[10034] = 8'b01100101;
DRAM[10035] = 8'b00100011;
DRAM[10036] = 8'b00100110;
DRAM[10037] = 8'b01000100;
DRAM[10038] = 8'b01001010;
DRAM[10039] = 8'b01001110;
DRAM[10040] = 8'b01101000;
DRAM[10041] = 8'b01111000;
DRAM[10042] = 8'b10000010;
DRAM[10043] = 8'b10000101;
DRAM[10044] = 8'b10001001;
DRAM[10045] = 8'b10001011;
DRAM[10046] = 8'b10010101;
DRAM[10047] = 8'b10010111;
DRAM[10048] = 8'b10011001;
DRAM[10049] = 8'b10011100;
DRAM[10050] = 8'b10100010;
DRAM[10051] = 8'b10100100;
DRAM[10052] = 8'b10100010;
DRAM[10053] = 8'b10011000;
DRAM[10054] = 8'b10010000;
DRAM[10055] = 8'b01111100;
DRAM[10056] = 8'b01111011;
DRAM[10057] = 8'b10000100;
DRAM[10058] = 8'b01111111;
DRAM[10059] = 8'b01111001;
DRAM[10060] = 8'b10000111;
DRAM[10061] = 8'b10100000;
DRAM[10062] = 8'b11001011;
DRAM[10063] = 8'b11011100;
DRAM[10064] = 8'b10010011;
DRAM[10065] = 8'b10010101;
DRAM[10066] = 8'b10010010;
DRAM[10067] = 8'b10000111;
DRAM[10068] = 8'b01111110;
DRAM[10069] = 8'b01100000;
DRAM[10070] = 8'b00101011;
DRAM[10071] = 8'b00110010;
DRAM[10072] = 8'b00111110;
DRAM[10073] = 8'b01000111;
DRAM[10074] = 8'b00111011;
DRAM[10075] = 8'b00101010;
DRAM[10076] = 8'b01111010;
DRAM[10077] = 8'b10011100;
DRAM[10078] = 8'b01101000;
DRAM[10079] = 8'b00101101;
DRAM[10080] = 8'b00101000;
DRAM[10081] = 8'b01100111;
DRAM[10082] = 8'b10001101;
DRAM[10083] = 8'b10010000;
DRAM[10084] = 8'b10100000;
DRAM[10085] = 8'b10011100;
DRAM[10086] = 8'b10011001;
DRAM[10087] = 8'b10011001;
DRAM[10088] = 8'b10010111;
DRAM[10089] = 8'b10010110;
DRAM[10090] = 8'b10010101;
DRAM[10091] = 8'b10010100;
DRAM[10092] = 8'b10010100;
DRAM[10093] = 8'b10010101;
DRAM[10094] = 8'b10010011;
DRAM[10095] = 8'b10001110;
DRAM[10096] = 8'b10001011;
DRAM[10097] = 8'b10001001;
DRAM[10098] = 8'b10000111;
DRAM[10099] = 8'b10101110;
DRAM[10100] = 8'b11000100;
DRAM[10101] = 8'b11000011;
DRAM[10102] = 8'b11000010;
DRAM[10103] = 8'b11000001;
DRAM[10104] = 8'b11001000;
DRAM[10105] = 8'b11010000;
DRAM[10106] = 8'b11010000;
DRAM[10107] = 8'b11001110;
DRAM[10108] = 8'b11001110;
DRAM[10109] = 8'b11001111;
DRAM[10110] = 8'b11010000;
DRAM[10111] = 8'b11001110;
DRAM[10112] = 8'b01010100;
DRAM[10113] = 8'b01010000;
DRAM[10114] = 8'b01001010;
DRAM[10115] = 8'b01000111;
DRAM[10116] = 8'b00111111;
DRAM[10117] = 8'b00110101;
DRAM[10118] = 8'b00110100;
DRAM[10119] = 8'b01110010;
DRAM[10120] = 8'b10010101;
DRAM[10121] = 8'b10101001;
DRAM[10122] = 8'b10101101;
DRAM[10123] = 8'b10110000;
DRAM[10124] = 8'b10110010;
DRAM[10125] = 8'b10101111;
DRAM[10126] = 8'b10011011;
DRAM[10127] = 8'b10000000;
DRAM[10128] = 8'b01010001;
DRAM[10129] = 8'b01011111;
DRAM[10130] = 8'b10000010;
DRAM[10131] = 8'b01101101;
DRAM[10132] = 8'b01101101;
DRAM[10133] = 8'b01110011;
DRAM[10134] = 8'b01000111;
DRAM[10135] = 8'b01001111;
DRAM[10136] = 8'b01100101;
DRAM[10137] = 8'b01011011;
DRAM[10138] = 8'b01001001;
DRAM[10139] = 8'b01000001;
DRAM[10140] = 8'b01101100;
DRAM[10141] = 8'b00111111;
DRAM[10142] = 8'b01100110;
DRAM[10143] = 8'b10001011;
DRAM[10144] = 8'b01000100;
DRAM[10145] = 8'b01011101;
DRAM[10146] = 8'b00111001;
DRAM[10147] = 8'b00110111;
DRAM[10148] = 8'b00110100;
DRAM[10149] = 8'b00101110;
DRAM[10150] = 8'b01000010;
DRAM[10151] = 8'b01010010;
DRAM[10152] = 8'b01000101;
DRAM[10153] = 8'b10000000;
DRAM[10154] = 8'b00111000;
DRAM[10155] = 8'b00100101;
DRAM[10156] = 8'b00100101;
DRAM[10157] = 8'b01001101;
DRAM[10158] = 8'b10100000;
DRAM[10159] = 8'b10001101;
DRAM[10160] = 8'b10001010;
DRAM[10161] = 8'b10100011;
DRAM[10162] = 8'b00111011;
DRAM[10163] = 8'b00100110;
DRAM[10164] = 8'b00101101;
DRAM[10165] = 8'b01000001;
DRAM[10166] = 8'b01010011;
DRAM[10167] = 8'b01001100;
DRAM[10168] = 8'b01101101;
DRAM[10169] = 8'b01111010;
DRAM[10170] = 8'b10000000;
DRAM[10171] = 8'b10000010;
DRAM[10172] = 8'b10000111;
DRAM[10173] = 8'b10001111;
DRAM[10174] = 8'b10010010;
DRAM[10175] = 8'b10010101;
DRAM[10176] = 8'b10011000;
DRAM[10177] = 8'b10011100;
DRAM[10178] = 8'b10011100;
DRAM[10179] = 8'b10011110;
DRAM[10180] = 8'b10011111;
DRAM[10181] = 8'b10010111;
DRAM[10182] = 8'b10001110;
DRAM[10183] = 8'b01110010;
DRAM[10184] = 8'b10000100;
DRAM[10185] = 8'b10001010;
DRAM[10186] = 8'b10001111;
DRAM[10187] = 8'b10000100;
DRAM[10188] = 8'b01111101;
DRAM[10189] = 8'b10011110;
DRAM[10190] = 8'b11001000;
DRAM[10191] = 8'b11011001;
DRAM[10192] = 8'b10001111;
DRAM[10193] = 8'b10010011;
DRAM[10194] = 8'b10001101;
DRAM[10195] = 8'b10000010;
DRAM[10196] = 8'b01110111;
DRAM[10197] = 8'b01000100;
DRAM[10198] = 8'b00101100;
DRAM[10199] = 8'b00110010;
DRAM[10200] = 8'b00111101;
DRAM[10201] = 8'b01000111;
DRAM[10202] = 8'b00111011;
DRAM[10203] = 8'b00101100;
DRAM[10204] = 8'b01011110;
DRAM[10205] = 8'b10011100;
DRAM[10206] = 8'b01111110;
DRAM[10207] = 8'b00101100;
DRAM[10208] = 8'b00101000;
DRAM[10209] = 8'b10000111;
DRAM[10210] = 8'b10010010;
DRAM[10211] = 8'b10010101;
DRAM[10212] = 8'b10011110;
DRAM[10213] = 8'b10011001;
DRAM[10214] = 8'b10011001;
DRAM[10215] = 8'b10010110;
DRAM[10216] = 8'b10010110;
DRAM[10217] = 8'b10010101;
DRAM[10218] = 8'b10010111;
DRAM[10219] = 8'b10010100;
DRAM[10220] = 8'b10010011;
DRAM[10221] = 8'b10010110;
DRAM[10222] = 8'b10010010;
DRAM[10223] = 8'b10010000;
DRAM[10224] = 8'b10001100;
DRAM[10225] = 8'b10000100;
DRAM[10226] = 8'b10010010;
DRAM[10227] = 8'b10111010;
DRAM[10228] = 8'b11000100;
DRAM[10229] = 8'b11000010;
DRAM[10230] = 8'b11000010;
DRAM[10231] = 8'b11000110;
DRAM[10232] = 8'b11001100;
DRAM[10233] = 8'b11001111;
DRAM[10234] = 8'b11001110;
DRAM[10235] = 8'b11001100;
DRAM[10236] = 8'b11001100;
DRAM[10237] = 8'b11010000;
DRAM[10238] = 8'b11010000;
DRAM[10239] = 8'b11001111;
DRAM[10240] = 8'b01010001;
DRAM[10241] = 8'b01010010;
DRAM[10242] = 8'b01001011;
DRAM[10243] = 8'b01001000;
DRAM[10244] = 8'b00111111;
DRAM[10245] = 8'b00111010;
DRAM[10246] = 8'b01000000;
DRAM[10247] = 8'b01110101;
DRAM[10248] = 8'b10010011;
DRAM[10249] = 8'b10100110;
DRAM[10250] = 8'b10101100;
DRAM[10251] = 8'b10101101;
DRAM[10252] = 8'b10110000;
DRAM[10253] = 8'b10101111;
DRAM[10254] = 8'b10011110;
DRAM[10255] = 8'b10000100;
DRAM[10256] = 8'b01100001;
DRAM[10257] = 8'b01011000;
DRAM[10258] = 8'b01011010;
DRAM[10259] = 8'b01100100;
DRAM[10260] = 8'b01101111;
DRAM[10261] = 8'b01101010;
DRAM[10262] = 8'b01001000;
DRAM[10263] = 8'b01010110;
DRAM[10264] = 8'b01110100;
DRAM[10265] = 8'b01011010;
DRAM[10266] = 8'b00110010;
DRAM[10267] = 8'b01110110;
DRAM[10268] = 8'b01001010;
DRAM[10269] = 8'b00110011;
DRAM[10270] = 8'b01101010;
DRAM[10271] = 8'b01111001;
DRAM[10272] = 8'b01101000;
DRAM[10273] = 8'b01101010;
DRAM[10274] = 8'b00101101;
DRAM[10275] = 8'b00110111;
DRAM[10276] = 8'b00111110;
DRAM[10277] = 8'b00100101;
DRAM[10278] = 8'b00110001;
DRAM[10279] = 8'b00110111;
DRAM[10280] = 8'b01010111;
DRAM[10281] = 8'b01011010;
DRAM[10282] = 8'b00101000;
DRAM[10283] = 8'b00101010;
DRAM[10284] = 8'b00100010;
DRAM[10285] = 8'b01101111;
DRAM[10286] = 8'b10110100;
DRAM[10287] = 8'b10110011;
DRAM[10288] = 8'b10111000;
DRAM[10289] = 8'b01001010;
DRAM[10290] = 8'b00100011;
DRAM[10291] = 8'b00101000;
DRAM[10292] = 8'b00101100;
DRAM[10293] = 8'b01000100;
DRAM[10294] = 8'b01010110;
DRAM[10295] = 8'b01010110;
DRAM[10296] = 8'b01101011;
DRAM[10297] = 8'b01111000;
DRAM[10298] = 8'b01111110;
DRAM[10299] = 8'b10000000;
DRAM[10300] = 8'b10001000;
DRAM[10301] = 8'b10001100;
DRAM[10302] = 8'b10010000;
DRAM[10303] = 8'b10010101;
DRAM[10304] = 8'b10011001;
DRAM[10305] = 8'b10011000;
DRAM[10306] = 8'b10011010;
DRAM[10307] = 8'b10011110;
DRAM[10308] = 8'b10011110;
DRAM[10309] = 8'b10011001;
DRAM[10310] = 8'b10010000;
DRAM[10311] = 8'b01110110;
DRAM[10312] = 8'b10000100;
DRAM[10313] = 8'b01100110;
DRAM[10314] = 8'b01011111;
DRAM[10315] = 8'b01110000;
DRAM[10316] = 8'b01111010;
DRAM[10317] = 8'b10001000;
DRAM[10318] = 8'b10111001;
DRAM[10319] = 8'b10111101;
DRAM[10320] = 8'b10010010;
DRAM[10321] = 8'b10010101;
DRAM[10322] = 8'b10001101;
DRAM[10323] = 8'b10000100;
DRAM[10324] = 8'b01101001;
DRAM[10325] = 8'b00101100;
DRAM[10326] = 8'b00101100;
DRAM[10327] = 8'b00110100;
DRAM[10328] = 8'b00111100;
DRAM[10329] = 8'b01000010;
DRAM[10330] = 8'b00110110;
DRAM[10331] = 8'b00101110;
DRAM[10332] = 8'b01011011;
DRAM[10333] = 8'b10100111;
DRAM[10334] = 8'b10000000;
DRAM[10335] = 8'b00101011;
DRAM[10336] = 8'b00111010;
DRAM[10337] = 8'b10001011;
DRAM[10338] = 8'b10001111;
DRAM[10339] = 8'b10011100;
DRAM[10340] = 8'b10011100;
DRAM[10341] = 8'b10011001;
DRAM[10342] = 8'b10011000;
DRAM[10343] = 8'b10010101;
DRAM[10344] = 8'b10010110;
DRAM[10345] = 8'b10010110;
DRAM[10346] = 8'b10010111;
DRAM[10347] = 8'b10010011;
DRAM[10348] = 8'b10010011;
DRAM[10349] = 8'b10010010;
DRAM[10350] = 8'b10010001;
DRAM[10351] = 8'b10001101;
DRAM[10352] = 8'b10001000;
DRAM[10353] = 8'b10000100;
DRAM[10354] = 8'b10100011;
DRAM[10355] = 8'b11000000;
DRAM[10356] = 8'b11000101;
DRAM[10357] = 8'b11000010;
DRAM[10358] = 8'b11000101;
DRAM[10359] = 8'b11001011;
DRAM[10360] = 8'b11001100;
DRAM[10361] = 8'b11001101;
DRAM[10362] = 8'b11001101;
DRAM[10363] = 8'b11001111;
DRAM[10364] = 8'b11010001;
DRAM[10365] = 8'b11010001;
DRAM[10366] = 8'b11010000;
DRAM[10367] = 8'b11001111;
DRAM[10368] = 8'b01001110;
DRAM[10369] = 8'b01001100;
DRAM[10370] = 8'b01001110;
DRAM[10371] = 8'b01001010;
DRAM[10372] = 8'b01000010;
DRAM[10373] = 8'b01000011;
DRAM[10374] = 8'b01010000;
DRAM[10375] = 8'b10000010;
DRAM[10376] = 8'b10011010;
DRAM[10377] = 8'b10100111;
DRAM[10378] = 8'b10101101;
DRAM[10379] = 8'b10101110;
DRAM[10380] = 8'b10110001;
DRAM[10381] = 8'b10110000;
DRAM[10382] = 8'b10011111;
DRAM[10383] = 8'b10000001;
DRAM[10384] = 8'b01010100;
DRAM[10385] = 8'b01001100;
DRAM[10386] = 8'b01011001;
DRAM[10387] = 8'b01100010;
DRAM[10388] = 8'b01101111;
DRAM[10389] = 8'b01100011;
DRAM[10390] = 8'b01010101;
DRAM[10391] = 8'b01011110;
DRAM[10392] = 8'b01100101;
DRAM[10393] = 8'b01000011;
DRAM[10394] = 8'b00111100;
DRAM[10395] = 8'b01110100;
DRAM[10396] = 8'b01001111;
DRAM[10397] = 8'b01000101;
DRAM[10398] = 8'b01110000;
DRAM[10399] = 8'b01100110;
DRAM[10400] = 8'b10000101;
DRAM[10401] = 8'b01101111;
DRAM[10402] = 8'b00011110;
DRAM[10403] = 8'b00110001;
DRAM[10404] = 8'b01001100;
DRAM[10405] = 8'b01000011;
DRAM[10406] = 8'b00100100;
DRAM[10407] = 8'b00101100;
DRAM[10408] = 8'b01110010;
DRAM[10409] = 8'b00110010;
DRAM[10410] = 8'b00110100;
DRAM[10411] = 8'b00111011;
DRAM[10412] = 8'b00111001;
DRAM[10413] = 8'b10001111;
DRAM[10414] = 8'b10100101;
DRAM[10415] = 8'b10110110;
DRAM[10416] = 8'b01010101;
DRAM[10417] = 8'b00100100;
DRAM[10418] = 8'b00101011;
DRAM[10419] = 8'b00101100;
DRAM[10420] = 8'b00101110;
DRAM[10421] = 8'b01001010;
DRAM[10422] = 8'b01100000;
DRAM[10423] = 8'b01011100;
DRAM[10424] = 8'b01101100;
DRAM[10425] = 8'b01111001;
DRAM[10426] = 8'b01111100;
DRAM[10427] = 8'b10000010;
DRAM[10428] = 8'b10000101;
DRAM[10429] = 8'b10001011;
DRAM[10430] = 8'b10010010;
DRAM[10431] = 8'b10010100;
DRAM[10432] = 8'b10010000;
DRAM[10433] = 8'b10010111;
DRAM[10434] = 8'b10011011;
DRAM[10435] = 8'b10011101;
DRAM[10436] = 8'b10011101;
DRAM[10437] = 8'b10011011;
DRAM[10438] = 8'b10010100;
DRAM[10439] = 8'b10000100;
DRAM[10440] = 8'b01111110;
DRAM[10441] = 8'b01110111;
DRAM[10442] = 8'b01111011;
DRAM[10443] = 8'b01110010;
DRAM[10444] = 8'b01101011;
DRAM[10445] = 8'b01111101;
DRAM[10446] = 8'b10110000;
DRAM[10447] = 8'b10101010;
DRAM[10448] = 8'b10011001;
DRAM[10449] = 8'b10001111;
DRAM[10450] = 8'b10001000;
DRAM[10451] = 8'b01111111;
DRAM[10452] = 8'b01001010;
DRAM[10453] = 8'b00110001;
DRAM[10454] = 8'b00101110;
DRAM[10455] = 8'b00111000;
DRAM[10456] = 8'b01000010;
DRAM[10457] = 8'b01000010;
DRAM[10458] = 8'b00110110;
DRAM[10459] = 8'b00101111;
DRAM[10460] = 8'b01001000;
DRAM[10461] = 8'b10100100;
DRAM[10462] = 8'b10000101;
DRAM[10463] = 8'b00111000;
DRAM[10464] = 8'b01100100;
DRAM[10465] = 8'b10010011;
DRAM[10466] = 8'b10010000;
DRAM[10467] = 8'b10011100;
DRAM[10468] = 8'b10011100;
DRAM[10469] = 8'b10011000;
DRAM[10470] = 8'b10010111;
DRAM[10471] = 8'b10010110;
DRAM[10472] = 8'b10010101;
DRAM[10473] = 8'b10010110;
DRAM[10474] = 8'b10010011;
DRAM[10475] = 8'b10010101;
DRAM[10476] = 8'b10010001;
DRAM[10477] = 8'b10010000;
DRAM[10478] = 8'b10010010;
DRAM[10479] = 8'b10001101;
DRAM[10480] = 8'b10001010;
DRAM[10481] = 8'b10000111;
DRAM[10482] = 8'b10101110;
DRAM[10483] = 8'b11000010;
DRAM[10484] = 8'b11000100;
DRAM[10485] = 8'b11000110;
DRAM[10486] = 8'b11001010;
DRAM[10487] = 8'b11001111;
DRAM[10488] = 8'b11010000;
DRAM[10489] = 8'b11001111;
DRAM[10490] = 8'b11001111;
DRAM[10491] = 8'b11010011;
DRAM[10492] = 8'b11010001;
DRAM[10493] = 8'b11010010;
DRAM[10494] = 8'b11010000;
DRAM[10495] = 8'b11001111;
DRAM[10496] = 8'b01010000;
DRAM[10497] = 8'b01001100;
DRAM[10498] = 8'b01001011;
DRAM[10499] = 8'b01001011;
DRAM[10500] = 8'b01000101;
DRAM[10501] = 8'b01001010;
DRAM[10502] = 8'b01011110;
DRAM[10503] = 8'b10000111;
DRAM[10504] = 8'b10011101;
DRAM[10505] = 8'b10100110;
DRAM[10506] = 8'b10101001;
DRAM[10507] = 8'b10101011;
DRAM[10508] = 8'b10110010;
DRAM[10509] = 8'b10110011;
DRAM[10510] = 8'b10011110;
DRAM[10511] = 8'b10000011;
DRAM[10512] = 8'b01010110;
DRAM[10513] = 8'b01001100;
DRAM[10514] = 8'b01011010;
DRAM[10515] = 8'b01100001;
DRAM[10516] = 8'b01110100;
DRAM[10517] = 8'b01110001;
DRAM[10518] = 8'b00101000;
DRAM[10519] = 8'b01010101;
DRAM[10520] = 8'b01000010;
DRAM[10521] = 8'b00110110;
DRAM[10522] = 8'b01101000;
DRAM[10523] = 8'b00111001;
DRAM[10524] = 8'b01001010;
DRAM[10525] = 8'b01001011;
DRAM[10526] = 8'b01101100;
DRAM[10527] = 8'b01101101;
DRAM[10528] = 8'b01110111;
DRAM[10529] = 8'b01110110;
DRAM[10530] = 8'b01000101;
DRAM[10531] = 8'b00101111;
DRAM[10532] = 8'b01010100;
DRAM[10533] = 8'b10010010;
DRAM[10534] = 8'b00100000;
DRAM[10535] = 8'b01000000;
DRAM[10536] = 8'b01001000;
DRAM[10537] = 8'b01000000;
DRAM[10538] = 8'b01100101;
DRAM[10539] = 8'b10000010;
DRAM[10540] = 8'b10010000;
DRAM[10541] = 8'b01101001;
DRAM[10542] = 8'b10001011;
DRAM[10543] = 8'b10100010;
DRAM[10544] = 8'b00101011;
DRAM[10545] = 8'b00101111;
DRAM[10546] = 8'b01000101;
DRAM[10547] = 8'b00110010;
DRAM[10548] = 8'b00101101;
DRAM[10549] = 8'b01001100;
DRAM[10550] = 8'b01101111;
DRAM[10551] = 8'b01011100;
DRAM[10552] = 8'b01110000;
DRAM[10553] = 8'b01111010;
DRAM[10554] = 8'b01111101;
DRAM[10555] = 8'b10000010;
DRAM[10556] = 8'b10000001;
DRAM[10557] = 8'b10001000;
DRAM[10558] = 8'b10010000;
DRAM[10559] = 8'b10010001;
DRAM[10560] = 8'b10010010;
DRAM[10561] = 8'b10010110;
DRAM[10562] = 8'b10011011;
DRAM[10563] = 8'b10011100;
DRAM[10564] = 8'b10011110;
DRAM[10565] = 8'b10011110;
DRAM[10566] = 8'b10011001;
DRAM[10567] = 8'b10010100;
DRAM[10568] = 8'b10001100;
DRAM[10569] = 8'b10000001;
DRAM[10570] = 8'b10001010;
DRAM[10571] = 8'b10001110;
DRAM[10572] = 8'b10010111;
DRAM[10573] = 8'b11000001;
DRAM[10574] = 8'b10111011;
DRAM[10575] = 8'b10100101;
DRAM[10576] = 8'b10010111;
DRAM[10577] = 8'b10001111;
DRAM[10578] = 8'b10000101;
DRAM[10579] = 8'b01110100;
DRAM[10580] = 8'b00110001;
DRAM[10581] = 8'b00101101;
DRAM[10582] = 8'b00110000;
DRAM[10583] = 8'b00111011;
DRAM[10584] = 8'b01001110;
DRAM[10585] = 8'b01001001;
DRAM[10586] = 8'b00110111;
DRAM[10587] = 8'b00111000;
DRAM[10588] = 8'b00110001;
DRAM[10589] = 8'b10100010;
DRAM[10590] = 8'b10000010;
DRAM[10591] = 8'b01001001;
DRAM[10592] = 8'b01110010;
DRAM[10593] = 8'b10010011;
DRAM[10594] = 8'b10010100;
DRAM[10595] = 8'b10011110;
DRAM[10596] = 8'b10011011;
DRAM[10597] = 8'b10011010;
DRAM[10598] = 8'b10010110;
DRAM[10599] = 8'b10010111;
DRAM[10600] = 8'b10010110;
DRAM[10601] = 8'b10010100;
DRAM[10602] = 8'b10010101;
DRAM[10603] = 8'b10010010;
DRAM[10604] = 8'b10010010;
DRAM[10605] = 8'b10001111;
DRAM[10606] = 8'b10001110;
DRAM[10607] = 8'b10001101;
DRAM[10608] = 8'b10000100;
DRAM[10609] = 8'b10010010;
DRAM[10610] = 8'b10111001;
DRAM[10611] = 8'b11000011;
DRAM[10612] = 8'b11000100;
DRAM[10613] = 8'b11001000;
DRAM[10614] = 8'b11001101;
DRAM[10615] = 8'b11010000;
DRAM[10616] = 8'b11001110;
DRAM[10617] = 8'b11001111;
DRAM[10618] = 8'b11010000;
DRAM[10619] = 8'b11010010;
DRAM[10620] = 8'b11010010;
DRAM[10621] = 8'b11010000;
DRAM[10622] = 8'b11010000;
DRAM[10623] = 8'b11010010;
DRAM[10624] = 8'b01010001;
DRAM[10625] = 8'b01001110;
DRAM[10626] = 8'b01001110;
DRAM[10627] = 8'b01001010;
DRAM[10628] = 8'b01000001;
DRAM[10629] = 8'b01000100;
DRAM[10630] = 8'b01100110;
DRAM[10631] = 8'b10001100;
DRAM[10632] = 8'b10011110;
DRAM[10633] = 8'b10100100;
DRAM[10634] = 8'b10101010;
DRAM[10635] = 8'b10101110;
DRAM[10636] = 8'b10110011;
DRAM[10637] = 8'b10110010;
DRAM[10638] = 8'b10100001;
DRAM[10639] = 8'b10000110;
DRAM[10640] = 8'b01011010;
DRAM[10641] = 8'b01001110;
DRAM[10642] = 8'b01011000;
DRAM[10643] = 8'b01100011;
DRAM[10644] = 8'b01111000;
DRAM[10645] = 8'b10001000;
DRAM[10646] = 8'b00110101;
DRAM[10647] = 8'b01001010;
DRAM[10648] = 8'b01010000;
DRAM[10649] = 8'b01101011;
DRAM[10650] = 8'b00111110;
DRAM[10651] = 8'b00110011;
DRAM[10652] = 8'b01001000;
DRAM[10653] = 8'b01010010;
DRAM[10654] = 8'b01011110;
DRAM[10655] = 8'b01110000;
DRAM[10656] = 8'b01101001;
DRAM[10657] = 8'b01111101;
DRAM[10658] = 8'b01101010;
DRAM[10659] = 8'b00111101;
DRAM[10660] = 8'b01010000;
DRAM[10661] = 8'b01010111;
DRAM[10662] = 8'b00111011;
DRAM[10663] = 8'b00101011;
DRAM[10664] = 8'b01001010;
DRAM[10665] = 8'b10000000;
DRAM[10666] = 8'b10010100;
DRAM[10667] = 8'b10110101;
DRAM[10668] = 8'b01010111;
DRAM[10669] = 8'b01110111;
DRAM[10670] = 8'b10101111;
DRAM[10671] = 8'b00101000;
DRAM[10672] = 8'b00110000;
DRAM[10673] = 8'b00110011;
DRAM[10674] = 8'b00111101;
DRAM[10675] = 8'b00111100;
DRAM[10676] = 8'b00110010;
DRAM[10677] = 8'b01001100;
DRAM[10678] = 8'b01110001;
DRAM[10679] = 8'b01011111;
DRAM[10680] = 8'b01110011;
DRAM[10681] = 8'b01111111;
DRAM[10682] = 8'b01111111;
DRAM[10683] = 8'b10000001;
DRAM[10684] = 8'b10000110;
DRAM[10685] = 8'b10001100;
DRAM[10686] = 8'b10001110;
DRAM[10687] = 8'b10001110;
DRAM[10688] = 8'b10001111;
DRAM[10689] = 8'b10010101;
DRAM[10690] = 8'b10011001;
DRAM[10691] = 8'b10011011;
DRAM[10692] = 8'b10011110;
DRAM[10693] = 8'b10011101;
DRAM[10694] = 8'b10011001;
DRAM[10695] = 8'b10010111;
DRAM[10696] = 8'b10010011;
DRAM[10697] = 8'b10010000;
DRAM[10698] = 8'b10100010;
DRAM[10699] = 8'b10111101;
DRAM[10700] = 8'b10101000;
DRAM[10701] = 8'b11000101;
DRAM[10702] = 8'b11000000;
DRAM[10703] = 8'b10100100;
DRAM[10704] = 8'b10010011;
DRAM[10705] = 8'b10001101;
DRAM[10706] = 8'b10000101;
DRAM[10707] = 8'b01001110;
DRAM[10708] = 8'b00110010;
DRAM[10709] = 8'b00101111;
DRAM[10710] = 8'b00110001;
DRAM[10711] = 8'b01000010;
DRAM[10712] = 8'b01010001;
DRAM[10713] = 8'b01000110;
DRAM[10714] = 8'b00111000;
DRAM[10715] = 8'b00111010;
DRAM[10716] = 8'b00101010;
DRAM[10717] = 8'b10100001;
DRAM[10718] = 8'b10000111;
DRAM[10719] = 8'b01010001;
DRAM[10720] = 8'b10000001;
DRAM[10721] = 8'b10010001;
DRAM[10722] = 8'b10010111;
DRAM[10723] = 8'b10011110;
DRAM[10724] = 8'b10011010;
DRAM[10725] = 8'b10011010;
DRAM[10726] = 8'b10010111;
DRAM[10727] = 8'b10010111;
DRAM[10728] = 8'b10010101;
DRAM[10729] = 8'b10010110;
DRAM[10730] = 8'b10010011;
DRAM[10731] = 8'b10010010;
DRAM[10732] = 8'b10010100;
DRAM[10733] = 8'b10010001;
DRAM[10734] = 8'b10001101;
DRAM[10735] = 8'b10001100;
DRAM[10736] = 8'b10000011;
DRAM[10737] = 8'b10010101;
DRAM[10738] = 8'b10111010;
DRAM[10739] = 8'b11000011;
DRAM[10740] = 8'b11000110;
DRAM[10741] = 8'b11001010;
DRAM[10742] = 8'b11010000;
DRAM[10743] = 8'b11001111;
DRAM[10744] = 8'b11001101;
DRAM[10745] = 8'b11001111;
DRAM[10746] = 8'b11010001;
DRAM[10747] = 8'b11010001;
DRAM[10748] = 8'b11010010;
DRAM[10749] = 8'b11010011;
DRAM[10750] = 8'b11010011;
DRAM[10751] = 8'b11010100;
DRAM[10752] = 8'b01001000;
DRAM[10753] = 8'b01001001;
DRAM[10754] = 8'b01001000;
DRAM[10755] = 8'b01000110;
DRAM[10756] = 8'b00111111;
DRAM[10757] = 8'b01000111;
DRAM[10758] = 8'b01101000;
DRAM[10759] = 8'b10001010;
DRAM[10760] = 8'b10011110;
DRAM[10761] = 8'b10100101;
DRAM[10762] = 8'b10101010;
DRAM[10763] = 8'b10101100;
DRAM[10764] = 8'b10110011;
DRAM[10765] = 8'b10110000;
DRAM[10766] = 8'b10100001;
DRAM[10767] = 8'b10000010;
DRAM[10768] = 8'b01010110;
DRAM[10769] = 8'b01001100;
DRAM[10770] = 8'b01010111;
DRAM[10771] = 8'b01101011;
DRAM[10772] = 8'b10001010;
DRAM[10773] = 8'b01101100;
DRAM[10774] = 8'b01000000;
DRAM[10775] = 8'b01010100;
DRAM[10776] = 8'b01111000;
DRAM[10777] = 8'b00110001;
DRAM[10778] = 8'b01000110;
DRAM[10779] = 8'b00110100;
DRAM[10780] = 8'b01001100;
DRAM[10781] = 8'b01000011;
DRAM[10782] = 8'b01001010;
DRAM[10783] = 8'b01101000;
DRAM[10784] = 8'b01001110;
DRAM[10785] = 8'b01110110;
DRAM[10786] = 8'b10001010;
DRAM[10787] = 8'b01000010;
DRAM[10788] = 8'b01101000;
DRAM[10789] = 8'b00111101;
DRAM[10790] = 8'b00101011;
DRAM[10791] = 8'b00111110;
DRAM[10792] = 8'b10000001;
DRAM[10793] = 8'b10011101;
DRAM[10794] = 8'b10110100;
DRAM[10795] = 8'b10000100;
DRAM[10796] = 8'b01011110;
DRAM[10797] = 8'b10010100;
DRAM[10798] = 8'b01001010;
DRAM[10799] = 8'b00101011;
DRAM[10800] = 8'b00110010;
DRAM[10801] = 8'b00110000;
DRAM[10802] = 8'b00110110;
DRAM[10803] = 8'b01000001;
DRAM[10804] = 8'b00101110;
DRAM[10805] = 8'b00111000;
DRAM[10806] = 8'b01100100;
DRAM[10807] = 8'b01011010;
DRAM[10808] = 8'b01110001;
DRAM[10809] = 8'b01111010;
DRAM[10810] = 8'b01111101;
DRAM[10811] = 8'b10000001;
DRAM[10812] = 8'b10000100;
DRAM[10813] = 8'b10001001;
DRAM[10814] = 8'b10001110;
DRAM[10815] = 8'b10001011;
DRAM[10816] = 8'b10001101;
DRAM[10817] = 8'b10001111;
DRAM[10818] = 8'b10010101;
DRAM[10819] = 8'b10011000;
DRAM[10820] = 8'b10010110;
DRAM[10821] = 8'b10011010;
DRAM[10822] = 8'b10010111;
DRAM[10823] = 8'b10010110;
DRAM[10824] = 8'b10010100;
DRAM[10825] = 8'b10011010;
DRAM[10826] = 8'b10110000;
DRAM[10827] = 8'b11001100;
DRAM[10828] = 8'b10110001;
DRAM[10829] = 8'b11001011;
DRAM[10830] = 8'b10111110;
DRAM[10831] = 8'b10100000;
DRAM[10832] = 8'b10010000;
DRAM[10833] = 8'b10001010;
DRAM[10834] = 8'b01111101;
DRAM[10835] = 8'b00101100;
DRAM[10836] = 8'b00110000;
DRAM[10837] = 8'b00101110;
DRAM[10838] = 8'b00110000;
DRAM[10839] = 8'b00111111;
DRAM[10840] = 8'b01010100;
DRAM[10841] = 8'b01000111;
DRAM[10842] = 8'b00111101;
DRAM[10843] = 8'b00110001;
DRAM[10844] = 8'b00101010;
DRAM[10845] = 8'b10010000;
DRAM[10846] = 8'b10000100;
DRAM[10847] = 8'b01100000;
DRAM[10848] = 8'b10001011;
DRAM[10849] = 8'b10010000;
DRAM[10850] = 8'b10011011;
DRAM[10851] = 8'b10011001;
DRAM[10852] = 8'b10011011;
DRAM[10853] = 8'b10010111;
DRAM[10854] = 8'b10010111;
DRAM[10855] = 8'b10010011;
DRAM[10856] = 8'b10010110;
DRAM[10857] = 8'b10010110;
DRAM[10858] = 8'b10010001;
DRAM[10859] = 8'b10010010;
DRAM[10860] = 8'b10010000;
DRAM[10861] = 8'b10001111;
DRAM[10862] = 8'b10001110;
DRAM[10863] = 8'b10001011;
DRAM[10864] = 8'b10000111;
DRAM[10865] = 8'b10011101;
DRAM[10866] = 8'b10111110;
DRAM[10867] = 8'b11000110;
DRAM[10868] = 8'b11000111;
DRAM[10869] = 8'b11010000;
DRAM[10870] = 8'b11010001;
DRAM[10871] = 8'b11001111;
DRAM[10872] = 8'b11010000;
DRAM[10873] = 8'b11001111;
DRAM[10874] = 8'b11010000;
DRAM[10875] = 8'b11010001;
DRAM[10876] = 8'b11010100;
DRAM[10877] = 8'b11010001;
DRAM[10878] = 8'b11010011;
DRAM[10879] = 8'b11010011;
DRAM[10880] = 8'b01000101;
DRAM[10881] = 8'b01000111;
DRAM[10882] = 8'b01000110;
DRAM[10883] = 8'b01000101;
DRAM[10884] = 8'b00111110;
DRAM[10885] = 8'b01001010;
DRAM[10886] = 8'b01100010;
DRAM[10887] = 8'b10000111;
DRAM[10888] = 8'b10011101;
DRAM[10889] = 8'b10100110;
DRAM[10890] = 8'b10101010;
DRAM[10891] = 8'b10101110;
DRAM[10892] = 8'b10110010;
DRAM[10893] = 8'b10110010;
DRAM[10894] = 8'b10100010;
DRAM[10895] = 8'b10000110;
DRAM[10896] = 8'b01010100;
DRAM[10897] = 8'b01001001;
DRAM[10898] = 8'b01011001;
DRAM[10899] = 8'b10000011;
DRAM[10900] = 8'b01101100;
DRAM[10901] = 8'b01101111;
DRAM[10902] = 8'b01001001;
DRAM[10903] = 8'b01100111;
DRAM[10904] = 8'b01001110;
DRAM[10905] = 8'b00110100;
DRAM[10906] = 8'b01000011;
DRAM[10907] = 8'b01000011;
DRAM[10908] = 8'b01000000;
DRAM[10909] = 8'b01010010;
DRAM[10910] = 8'b01000010;
DRAM[10911] = 8'b01011010;
DRAM[10912] = 8'b01000010;
DRAM[10913] = 8'b01101111;
DRAM[10914] = 8'b01110111;
DRAM[10915] = 8'b10001011;
DRAM[10916] = 8'b01000001;
DRAM[10917] = 8'b00101011;
DRAM[10918] = 8'b01100011;
DRAM[10919] = 8'b01101101;
DRAM[10920] = 8'b01111001;
DRAM[10921] = 8'b10101001;
DRAM[10922] = 8'b10100001;
DRAM[10923] = 8'b01011111;
DRAM[10924] = 8'b01110110;
DRAM[10925] = 8'b01011100;
DRAM[10926] = 8'b00100111;
DRAM[10927] = 8'b00111101;
DRAM[10928] = 8'b00110011;
DRAM[10929] = 8'b00101111;
DRAM[10930] = 8'b00110011;
DRAM[10931] = 8'b01000111;
DRAM[10932] = 8'b00110010;
DRAM[10933] = 8'b00110000;
DRAM[10934] = 8'b01100010;
DRAM[10935] = 8'b01011100;
DRAM[10936] = 8'b01101101;
DRAM[10937] = 8'b01110111;
DRAM[10938] = 8'b01111101;
DRAM[10939] = 8'b10000000;
DRAM[10940] = 8'b10000111;
DRAM[10941] = 8'b10001011;
DRAM[10942] = 8'b10001110;
DRAM[10943] = 8'b10001110;
DRAM[10944] = 8'b10001010;
DRAM[10945] = 8'b10001101;
DRAM[10946] = 8'b10001101;
DRAM[10947] = 8'b10010001;
DRAM[10948] = 8'b10010010;
DRAM[10949] = 8'b10010100;
DRAM[10950] = 8'b10010010;
DRAM[10951] = 8'b10010010;
DRAM[10952] = 8'b10011000;
DRAM[10953] = 8'b10011111;
DRAM[10954] = 8'b10110111;
DRAM[10955] = 8'b11001111;
DRAM[10956] = 8'b10111001;
DRAM[10957] = 8'b11001010;
DRAM[10958] = 8'b11000000;
DRAM[10959] = 8'b10011011;
DRAM[10960] = 8'b10001100;
DRAM[10961] = 8'b10001010;
DRAM[10962] = 8'b01011010;
DRAM[10963] = 8'b00101100;
DRAM[10964] = 8'b00110100;
DRAM[10965] = 8'b00101110;
DRAM[10966] = 8'b00110100;
DRAM[10967] = 8'b01000100;
DRAM[10968] = 8'b01010010;
DRAM[10969] = 8'b01000110;
DRAM[10970] = 8'b00111001;
DRAM[10971] = 8'b00110110;
DRAM[10972] = 8'b00101000;
DRAM[10973] = 8'b10001010;
DRAM[10974] = 8'b10001111;
DRAM[10975] = 8'b01100110;
DRAM[10976] = 8'b10001011;
DRAM[10977] = 8'b10010000;
DRAM[10978] = 8'b10011011;
DRAM[10979] = 8'b10011010;
DRAM[10980] = 8'b10011000;
DRAM[10981] = 8'b10011000;
DRAM[10982] = 8'b10010100;
DRAM[10983] = 8'b10010011;
DRAM[10984] = 8'b10010010;
DRAM[10985] = 8'b10010100;
DRAM[10986] = 8'b10010101;
DRAM[10987] = 8'b10010010;
DRAM[10988] = 8'b10010001;
DRAM[10989] = 8'b10010001;
DRAM[10990] = 8'b10001101;
DRAM[10991] = 8'b10000110;
DRAM[10992] = 8'b10000000;
DRAM[10993] = 8'b10100010;
DRAM[10994] = 8'b11000001;
DRAM[10995] = 8'b11000111;
DRAM[10996] = 8'b11001101;
DRAM[10997] = 8'b11010000;
DRAM[10998] = 8'b11010000;
DRAM[10999] = 8'b11010000;
DRAM[11000] = 8'b11010000;
DRAM[11001] = 8'b11001111;
DRAM[11002] = 8'b11001111;
DRAM[11003] = 8'b11010010;
DRAM[11004] = 8'b11010011;
DRAM[11005] = 8'b11010011;
DRAM[11006] = 8'b11010101;
DRAM[11007] = 8'b11010011;
DRAM[11008] = 8'b01000010;
DRAM[11009] = 8'b00111111;
DRAM[11010] = 8'b01000011;
DRAM[11011] = 8'b01000011;
DRAM[11012] = 8'b00111111;
DRAM[11013] = 8'b01000110;
DRAM[11014] = 8'b01100000;
DRAM[11015] = 8'b10001010;
DRAM[11016] = 8'b10011110;
DRAM[11017] = 8'b10101000;
DRAM[11018] = 8'b10101100;
DRAM[11019] = 8'b10101111;
DRAM[11020] = 8'b10110100;
DRAM[11021] = 8'b10110011;
DRAM[11022] = 8'b10100010;
DRAM[11023] = 8'b10000011;
DRAM[11024] = 8'b01010110;
DRAM[11025] = 8'b01001011;
DRAM[11026] = 8'b01111000;
DRAM[11027] = 8'b01011111;
DRAM[11028] = 8'b01101010;
DRAM[11029] = 8'b01100000;
DRAM[11030] = 8'b00110101;
DRAM[11031] = 8'b01010101;
DRAM[11032] = 8'b01001010;
DRAM[11033] = 8'b00111111;
DRAM[11034] = 8'b00111111;
DRAM[11035] = 8'b00111110;
DRAM[11036] = 8'b01011000;
DRAM[11037] = 8'b01011001;
DRAM[11038] = 8'b01010110;
DRAM[11039] = 8'b01010000;
DRAM[11040] = 8'b01011001;
DRAM[11041] = 8'b00111110;
DRAM[11042] = 8'b01100100;
DRAM[11043] = 8'b10000110;
DRAM[11044] = 8'b00111111;
DRAM[11045] = 8'b01010000;
DRAM[11046] = 8'b10000011;
DRAM[11047] = 8'b10111011;
DRAM[11048] = 8'b10111011;
DRAM[11049] = 8'b10110110;
DRAM[11050] = 8'b01100010;
DRAM[11051] = 8'b01100101;
DRAM[11052] = 8'b10001101;
DRAM[11053] = 8'b00101000;
DRAM[11054] = 8'b00101000;
DRAM[11055] = 8'b01010000;
DRAM[11056] = 8'b00110000;
DRAM[11057] = 8'b00101111;
DRAM[11058] = 8'b00111100;
DRAM[11059] = 8'b01001010;
DRAM[11060] = 8'b00101111;
DRAM[11061] = 8'b00110011;
DRAM[11062] = 8'b01100010;
DRAM[11063] = 8'b01010110;
DRAM[11064] = 8'b01100011;
DRAM[11065] = 8'b01110101;
DRAM[11066] = 8'b01111111;
DRAM[11067] = 8'b10000010;
DRAM[11068] = 8'b10000001;
DRAM[11069] = 8'b10001001;
DRAM[11070] = 8'b10001010;
DRAM[11071] = 8'b10001101;
DRAM[11072] = 8'b10001001;
DRAM[11073] = 8'b10001011;
DRAM[11074] = 8'b10000111;
DRAM[11075] = 8'b10000100;
DRAM[11076] = 8'b10001000;
DRAM[11077] = 8'b10001101;
DRAM[11078] = 8'b10001101;
DRAM[11079] = 8'b10001100;
DRAM[11080] = 8'b10010000;
DRAM[11081] = 8'b10001110;
DRAM[11082] = 8'b10001001;
DRAM[11083] = 8'b10010110;
DRAM[11084] = 8'b10100101;
DRAM[11085] = 8'b10010101;
DRAM[11086] = 8'b10011000;
DRAM[11087] = 8'b01111100;
DRAM[11088] = 8'b10000110;
DRAM[11089] = 8'b10001000;
DRAM[11090] = 8'b00101111;
DRAM[11091] = 8'b00101101;
DRAM[11092] = 8'b00110011;
DRAM[11093] = 8'b00110001;
DRAM[11094] = 8'b00111000;
DRAM[11095] = 8'b01000101;
DRAM[11096] = 8'b01010111;
DRAM[11097] = 8'b01001111;
DRAM[11098] = 8'b00111101;
DRAM[11099] = 8'b00111010;
DRAM[11100] = 8'b00101000;
DRAM[11101] = 8'b01110000;
DRAM[11102] = 8'b10001111;
DRAM[11103] = 8'b01110110;
DRAM[11104] = 8'b10001111;
DRAM[11105] = 8'b10001111;
DRAM[11106] = 8'b10011100;
DRAM[11107] = 8'b10011011;
DRAM[11108] = 8'b10011010;
DRAM[11109] = 8'b10010101;
DRAM[11110] = 8'b10010101;
DRAM[11111] = 8'b10010010;
DRAM[11112] = 8'b10010111;
DRAM[11113] = 8'b10010011;
DRAM[11114] = 8'b10010001;
DRAM[11115] = 8'b10010000;
DRAM[11116] = 8'b10010001;
DRAM[11117] = 8'b10001111;
DRAM[11118] = 8'b10001011;
DRAM[11119] = 8'b10001001;
DRAM[11120] = 8'b10000001;
DRAM[11121] = 8'b10100110;
DRAM[11122] = 8'b11000001;
DRAM[11123] = 8'b11001011;
DRAM[11124] = 8'b11010001;
DRAM[11125] = 8'b11010001;
DRAM[11126] = 8'b11010000;
DRAM[11127] = 8'b11010001;
DRAM[11128] = 8'b11010001;
DRAM[11129] = 8'b11010001;
DRAM[11130] = 8'b11010010;
DRAM[11131] = 8'b11010101;
DRAM[11132] = 8'b11010101;
DRAM[11133] = 8'b11010100;
DRAM[11134] = 8'b11010101;
DRAM[11135] = 8'b11010100;
DRAM[11136] = 8'b00111000;
DRAM[11137] = 8'b00111011;
DRAM[11138] = 8'b00111111;
DRAM[11139] = 8'b01000001;
DRAM[11140] = 8'b00111111;
DRAM[11141] = 8'b01001010;
DRAM[11142] = 8'b01100100;
DRAM[11143] = 8'b10001100;
DRAM[11144] = 8'b10011110;
DRAM[11145] = 8'b10101010;
DRAM[11146] = 8'b10101111;
DRAM[11147] = 8'b10110010;
DRAM[11148] = 8'b10110010;
DRAM[11149] = 8'b10110010;
DRAM[11150] = 8'b10100000;
DRAM[11151] = 8'b10000000;
DRAM[11152] = 8'b01010011;
DRAM[11153] = 8'b01100100;
DRAM[11154] = 8'b01101010;
DRAM[11155] = 8'b01011011;
DRAM[11156] = 8'b10001110;
DRAM[11157] = 8'b01011100;
DRAM[11158] = 8'b00111010;
DRAM[11159] = 8'b00111010;
DRAM[11160] = 8'b01000000;
DRAM[11161] = 8'b00111110;
DRAM[11162] = 8'b01000010;
DRAM[11163] = 8'b00111010;
DRAM[11164] = 8'b01010110;
DRAM[11165] = 8'b01110010;
DRAM[11166] = 8'b01101000;
DRAM[11167] = 8'b01011001;
DRAM[11168] = 8'b01000101;
DRAM[11169] = 8'b01100110;
DRAM[11170] = 8'b01011110;
DRAM[11171] = 8'b01010100;
DRAM[11172] = 8'b01010101;
DRAM[11173] = 8'b10001110;
DRAM[11174] = 8'b10001011;
DRAM[11175] = 8'b11000111;
DRAM[11176] = 8'b11001100;
DRAM[11177] = 8'b01101110;
DRAM[11178] = 8'b01100001;
DRAM[11179] = 8'b10100000;
DRAM[11180] = 8'b00111000;
DRAM[11181] = 8'b00101110;
DRAM[11182] = 8'b00101011;
DRAM[11183] = 8'b01000010;
DRAM[11184] = 8'b00101011;
DRAM[11185] = 8'b00110001;
DRAM[11186] = 8'b00111110;
DRAM[11187] = 8'b01001000;
DRAM[11188] = 8'b00111010;
DRAM[11189] = 8'b00101011;
DRAM[11190] = 8'b01100100;
DRAM[11191] = 8'b01011001;
DRAM[11192] = 8'b01011100;
DRAM[11193] = 8'b01110001;
DRAM[11194] = 8'b01111110;
DRAM[11195] = 8'b01111110;
DRAM[11196] = 8'b10000010;
DRAM[11197] = 8'b10000010;
DRAM[11198] = 8'b10001000;
DRAM[11199] = 8'b10010001;
DRAM[11200] = 8'b10010000;
DRAM[11201] = 8'b10010000;
DRAM[11202] = 8'b01100010;
DRAM[11203] = 8'b01011010;
DRAM[11204] = 8'b01100110;
DRAM[11205] = 8'b01101011;
DRAM[11206] = 8'b01101100;
DRAM[11207] = 8'b01110001;
DRAM[11208] = 8'b01101010;
DRAM[11209] = 8'b01100001;
DRAM[11210] = 8'b01101010;
DRAM[11211] = 8'b01111000;
DRAM[11212] = 8'b01110110;
DRAM[11213] = 8'b01011100;
DRAM[11214] = 8'b01110000;
DRAM[11215] = 8'b01110110;
DRAM[11216] = 8'b10001111;
DRAM[11217] = 8'b01011101;
DRAM[11218] = 8'b00101100;
DRAM[11219] = 8'b00110001;
DRAM[11220] = 8'b00110001;
DRAM[11221] = 8'b00110011;
DRAM[11222] = 8'b00111100;
DRAM[11223] = 8'b00111111;
DRAM[11224] = 8'b01010010;
DRAM[11225] = 8'b01001110;
DRAM[11226] = 8'b00110111;
DRAM[11227] = 8'b01000100;
DRAM[11228] = 8'b00101000;
DRAM[11229] = 8'b01100000;
DRAM[11230] = 8'b10001100;
DRAM[11231] = 8'b10001011;
DRAM[11232] = 8'b10010010;
DRAM[11233] = 8'b10010011;
DRAM[11234] = 8'b10011011;
DRAM[11235] = 8'b10011011;
DRAM[11236] = 8'b10010111;
DRAM[11237] = 8'b10011001;
DRAM[11238] = 8'b10010101;
DRAM[11239] = 8'b10010011;
DRAM[11240] = 8'b10010110;
DRAM[11241] = 8'b10010010;
DRAM[11242] = 8'b10010100;
DRAM[11243] = 8'b10010000;
DRAM[11244] = 8'b10010001;
DRAM[11245] = 8'b10001111;
DRAM[11246] = 8'b10001101;
DRAM[11247] = 8'b10000101;
DRAM[11248] = 8'b10000010;
DRAM[11249] = 8'b10101001;
DRAM[11250] = 8'b11000101;
DRAM[11251] = 8'b11010000;
DRAM[11252] = 8'b11010011;
DRAM[11253] = 8'b11010010;
DRAM[11254] = 8'b11010010;
DRAM[11255] = 8'b11010000;
DRAM[11256] = 8'b11010001;
DRAM[11257] = 8'b11010001;
DRAM[11258] = 8'b11010011;
DRAM[11259] = 8'b11010100;
DRAM[11260] = 8'b11010101;
DRAM[11261] = 8'b11010110;
DRAM[11262] = 8'b11010100;
DRAM[11263] = 8'b11010101;
DRAM[11264] = 8'b00111000;
DRAM[11265] = 8'b00111010;
DRAM[11266] = 8'b00111100;
DRAM[11267] = 8'b00111111;
DRAM[11268] = 8'b01000001;
DRAM[11269] = 8'b01010000;
DRAM[11270] = 8'b01100111;
DRAM[11271] = 8'b10001101;
DRAM[11272] = 8'b10100000;
DRAM[11273] = 8'b10101011;
DRAM[11274] = 8'b10110000;
DRAM[11275] = 8'b10110000;
DRAM[11276] = 8'b10110110;
DRAM[11277] = 8'b10110001;
DRAM[11278] = 8'b10100000;
DRAM[11279] = 8'b10000010;
DRAM[11280] = 8'b01101110;
DRAM[11281] = 8'b01111000;
DRAM[11282] = 8'b01010010;
DRAM[11283] = 8'b01111000;
DRAM[11284] = 8'b01111111;
DRAM[11285] = 8'b01010110;
DRAM[11286] = 8'b00111100;
DRAM[11287] = 8'b00111100;
DRAM[11288] = 8'b00110000;
DRAM[11289] = 8'b00110100;
DRAM[11290] = 8'b01001000;
DRAM[11291] = 8'b01000111;
DRAM[11292] = 8'b01100001;
DRAM[11293] = 8'b01111011;
DRAM[11294] = 8'b01010100;
DRAM[11295] = 8'b01100100;
DRAM[11296] = 8'b01100100;
DRAM[11297] = 8'b01011100;
DRAM[11298] = 8'b01100011;
DRAM[11299] = 8'b01010100;
DRAM[11300] = 8'b01110000;
DRAM[11301] = 8'b10010001;
DRAM[11302] = 8'b01111100;
DRAM[11303] = 8'b11010100;
DRAM[11304] = 8'b10011010;
DRAM[11305] = 8'b01100011;
DRAM[11306] = 8'b10001110;
DRAM[11307] = 8'b01100110;
DRAM[11308] = 8'b00101111;
DRAM[11309] = 8'b00110100;
DRAM[11310] = 8'b00101001;
DRAM[11311] = 8'b00111000;
DRAM[11312] = 8'b00110010;
DRAM[11313] = 8'b00110101;
DRAM[11314] = 8'b00111011;
DRAM[11315] = 8'b00111011;
DRAM[11316] = 8'b00111110;
DRAM[11317] = 8'b00110001;
DRAM[11318] = 8'b01011010;
DRAM[11319] = 8'b01010000;
DRAM[11320] = 8'b01011000;
DRAM[11321] = 8'b01101100;
DRAM[11322] = 8'b01111000;
DRAM[11323] = 8'b01111101;
DRAM[11324] = 8'b01111100;
DRAM[11325] = 8'b10000000;
DRAM[11326] = 8'b10001000;
DRAM[11327] = 8'b10001010;
DRAM[11328] = 8'b10010010;
DRAM[11329] = 8'b10010000;
DRAM[11330] = 8'b10000111;
DRAM[11331] = 8'b01111111;
DRAM[11332] = 8'b01111000;
DRAM[11333] = 8'b01110110;
DRAM[11334] = 8'b01111010;
DRAM[11335] = 8'b10000010;
DRAM[11336] = 8'b10001011;
DRAM[11337] = 8'b10011000;
DRAM[11338] = 8'b10010111;
DRAM[11339] = 8'b10101100;
DRAM[11340] = 8'b10101011;
DRAM[11341] = 8'b10001000;
DRAM[11342] = 8'b10001100;
DRAM[11343] = 8'b10010000;
DRAM[11344] = 8'b10000011;
DRAM[11345] = 8'b00101010;
DRAM[11346] = 8'b00101101;
DRAM[11347] = 8'b00110100;
DRAM[11348] = 8'b00101110;
DRAM[11349] = 8'b00110110;
DRAM[11350] = 8'b00111011;
DRAM[11351] = 8'b00111111;
DRAM[11352] = 8'b01001010;
DRAM[11353] = 8'b01001101;
DRAM[11354] = 8'b00111010;
DRAM[11355] = 8'b01001101;
DRAM[11356] = 8'b00101011;
DRAM[11357] = 8'b01010001;
DRAM[11358] = 8'b10010001;
DRAM[11359] = 8'b10011000;
DRAM[11360] = 8'b10010110;
DRAM[11361] = 8'b10010101;
DRAM[11362] = 8'b10011011;
DRAM[11363] = 8'b10011010;
DRAM[11364] = 8'b10011000;
DRAM[11365] = 8'b10011001;
DRAM[11366] = 8'b10011000;
DRAM[11367] = 8'b10010110;
DRAM[11368] = 8'b10010011;
DRAM[11369] = 8'b10010011;
DRAM[11370] = 8'b10010100;
DRAM[11371] = 8'b10010001;
DRAM[11372] = 8'b10010010;
DRAM[11373] = 8'b10010000;
DRAM[11374] = 8'b10001011;
DRAM[11375] = 8'b10000101;
DRAM[11376] = 8'b10000010;
DRAM[11377] = 8'b10110011;
DRAM[11378] = 8'b11001011;
DRAM[11379] = 8'b11010011;
DRAM[11380] = 8'b11010011;
DRAM[11381] = 8'b11010001;
DRAM[11382] = 8'b11010011;
DRAM[11383] = 8'b11010010;
DRAM[11384] = 8'b11010010;
DRAM[11385] = 8'b11010011;
DRAM[11386] = 8'b11010100;
DRAM[11387] = 8'b11010101;
DRAM[11388] = 8'b11010101;
DRAM[11389] = 8'b11010101;
DRAM[11390] = 8'b11010100;
DRAM[11391] = 8'b11010100;
DRAM[11392] = 8'b00110111;
DRAM[11393] = 8'b00111000;
DRAM[11394] = 8'b00111111;
DRAM[11395] = 8'b00111101;
DRAM[11396] = 8'b00111001;
DRAM[11397] = 8'b01010011;
DRAM[11398] = 8'b01100110;
DRAM[11399] = 8'b10001010;
DRAM[11400] = 8'b10011110;
DRAM[11401] = 8'b10101010;
DRAM[11402] = 8'b10110000;
DRAM[11403] = 8'b10110011;
DRAM[11404] = 8'b10110101;
DRAM[11405] = 8'b10110000;
DRAM[11406] = 8'b10100111;
DRAM[11407] = 8'b10001011;
DRAM[11408] = 8'b01111000;
DRAM[11409] = 8'b01000100;
DRAM[11410] = 8'b01011000;
DRAM[11411] = 8'b10001010;
DRAM[11412] = 8'b01101011;
DRAM[11413] = 8'b01001110;
DRAM[11414] = 8'b01001100;
DRAM[11415] = 8'b01011111;
DRAM[11416] = 8'b00101010;
DRAM[11417] = 8'b00110110;
DRAM[11418] = 8'b01010111;
DRAM[11419] = 8'b01010010;
DRAM[11420] = 8'b01101001;
DRAM[11421] = 8'b10000110;
DRAM[11422] = 8'b01000000;
DRAM[11423] = 8'b01011000;
DRAM[11424] = 8'b01100111;
DRAM[11425] = 8'b01011001;
DRAM[11426] = 8'b01001010;
DRAM[11427] = 8'b01100101;
DRAM[11428] = 8'b10000010;
DRAM[11429] = 8'b10010100;
DRAM[11430] = 8'b10000100;
DRAM[11431] = 8'b10110101;
DRAM[11432] = 8'b01101001;
DRAM[11433] = 8'b10010011;
DRAM[11434] = 8'b10010101;
DRAM[11435] = 8'b00101111;
DRAM[11436] = 8'b00110011;
DRAM[11437] = 8'b00110101;
DRAM[11438] = 8'b00101101;
DRAM[11439] = 8'b00110001;
DRAM[11440] = 8'b00110011;
DRAM[11441] = 8'b00110000;
DRAM[11442] = 8'b00111010;
DRAM[11443] = 8'b00111100;
DRAM[11444] = 8'b01000100;
DRAM[11445] = 8'b00110010;
DRAM[11446] = 8'b01000010;
DRAM[11447] = 8'b01001111;
DRAM[11448] = 8'b01001100;
DRAM[11449] = 8'b01100110;
DRAM[11450] = 8'b01101110;
DRAM[11451] = 8'b01110110;
DRAM[11452] = 8'b01111000;
DRAM[11453] = 8'b01111100;
DRAM[11454] = 8'b10000000;
DRAM[11455] = 8'b10000101;
DRAM[11456] = 8'b10010001;
DRAM[11457] = 8'b10010001;
DRAM[11458] = 8'b10001111;
DRAM[11459] = 8'b10000110;
DRAM[11460] = 8'b01111110;
DRAM[11461] = 8'b01111111;
DRAM[11462] = 8'b01111110;
DRAM[11463] = 8'b10000000;
DRAM[11464] = 8'b10010011;
DRAM[11465] = 8'b10011111;
DRAM[11466] = 8'b10100010;
DRAM[11467] = 8'b10011110;
DRAM[11468] = 8'b10100101;
DRAM[11469] = 8'b10001010;
DRAM[11470] = 8'b10010011;
DRAM[11471] = 8'b10001110;
DRAM[11472] = 8'b01010000;
DRAM[11473] = 8'b00101101;
DRAM[11474] = 8'b00101111;
DRAM[11475] = 8'b00110010;
DRAM[11476] = 8'b00101010;
DRAM[11477] = 8'b00111000;
DRAM[11478] = 8'b00110111;
DRAM[11479] = 8'b01000010;
DRAM[11480] = 8'b01001110;
DRAM[11481] = 8'b01001110;
DRAM[11482] = 8'b00111111;
DRAM[11483] = 8'b01001001;
DRAM[11484] = 8'b00101110;
DRAM[11485] = 8'b01000101;
DRAM[11486] = 8'b10011100;
DRAM[11487] = 8'b10010101;
DRAM[11488] = 8'b10010110;
DRAM[11489] = 8'b10011000;
DRAM[11490] = 8'b10011100;
DRAM[11491] = 8'b10011100;
DRAM[11492] = 8'b10011011;
DRAM[11493] = 8'b10010111;
DRAM[11494] = 8'b10011000;
DRAM[11495] = 8'b10011000;
DRAM[11496] = 8'b10010101;
DRAM[11497] = 8'b10010100;
DRAM[11498] = 8'b10010010;
DRAM[11499] = 8'b10001111;
DRAM[11500] = 8'b10010010;
DRAM[11501] = 8'b10010000;
DRAM[11502] = 8'b10001100;
DRAM[11503] = 8'b10000011;
DRAM[11504] = 8'b10000011;
DRAM[11505] = 8'b10110111;
DRAM[11506] = 8'b11001111;
DRAM[11507] = 8'b11010110;
DRAM[11508] = 8'b11010100;
DRAM[11509] = 8'b11010011;
DRAM[11510] = 8'b11010100;
DRAM[11511] = 8'b11010100;
DRAM[11512] = 8'b11010101;
DRAM[11513] = 8'b11010100;
DRAM[11514] = 8'b11010110;
DRAM[11515] = 8'b11010101;
DRAM[11516] = 8'b11010010;
DRAM[11517] = 8'b11010001;
DRAM[11518] = 8'b11010000;
DRAM[11519] = 8'b11001111;
DRAM[11520] = 8'b00110011;
DRAM[11521] = 8'b00110101;
DRAM[11522] = 8'b00110111;
DRAM[11523] = 8'b00111000;
DRAM[11524] = 8'b00111001;
DRAM[11525] = 8'b01010100;
DRAM[11526] = 8'b01100000;
DRAM[11527] = 8'b10001000;
DRAM[11528] = 8'b10011100;
DRAM[11529] = 8'b10101000;
DRAM[11530] = 8'b10110001;
DRAM[11531] = 8'b10110010;
DRAM[11532] = 8'b10110010;
DRAM[11533] = 8'b10110001;
DRAM[11534] = 8'b10100010;
DRAM[11535] = 8'b10000111;
DRAM[11536] = 8'b01010000;
DRAM[11537] = 8'b01001000;
DRAM[11538] = 8'b01111100;
DRAM[11539] = 8'b01110101;
DRAM[11540] = 8'b01101111;
DRAM[11541] = 8'b00111110;
DRAM[11542] = 8'b01101011;
DRAM[11543] = 8'b00111100;
DRAM[11544] = 8'b00101111;
DRAM[11545] = 8'b01000111;
DRAM[11546] = 8'b01000010;
DRAM[11547] = 8'b01011100;
DRAM[11548] = 8'b01111100;
DRAM[11549] = 8'b01011111;
DRAM[11550] = 8'b01100111;
DRAM[11551] = 8'b01100111;
DRAM[11552] = 8'b01000100;
DRAM[11553] = 8'b01110100;
DRAM[11554] = 8'b01100011;
DRAM[11555] = 8'b01101100;
DRAM[11556] = 8'b10011111;
DRAM[11557] = 8'b10001001;
DRAM[11558] = 8'b10010000;
DRAM[11559] = 8'b10011110;
DRAM[11560] = 8'b10011010;
DRAM[11561] = 8'b10100000;
DRAM[11562] = 8'b00111010;
DRAM[11563] = 8'b00111000;
DRAM[11564] = 8'b00110111;
DRAM[11565] = 8'b00111011;
DRAM[11566] = 8'b00110110;
DRAM[11567] = 8'b00110101;
DRAM[11568] = 8'b00110010;
DRAM[11569] = 8'b00111001;
DRAM[11570] = 8'b00111100;
DRAM[11571] = 8'b00111110;
DRAM[11572] = 8'b01000101;
DRAM[11573] = 8'b00110101;
DRAM[11574] = 8'b01000101;
DRAM[11575] = 8'b01010000;
DRAM[11576] = 8'b01000110;
DRAM[11577] = 8'b01011100;
DRAM[11578] = 8'b01101001;
DRAM[11579] = 8'b01101111;
DRAM[11580] = 8'b01110110;
DRAM[11581] = 8'b01110111;
DRAM[11582] = 8'b10000000;
DRAM[11583] = 8'b10000011;
DRAM[11584] = 8'b10001010;
DRAM[11585] = 8'b10001101;
DRAM[11586] = 8'b10001111;
DRAM[11587] = 8'b10001001;
DRAM[11588] = 8'b10000100;
DRAM[11589] = 8'b01111110;
DRAM[11590] = 8'b01111110;
DRAM[11591] = 8'b01111011;
DRAM[11592] = 8'b10000000;
DRAM[11593] = 8'b10000110;
DRAM[11594] = 8'b10001010;
DRAM[11595] = 8'b10000101;
DRAM[11596] = 8'b10001000;
DRAM[11597] = 8'b10010011;
DRAM[11598] = 8'b10010010;
DRAM[11599] = 8'b01110110;
DRAM[11600] = 8'b00110001;
DRAM[11601] = 8'b00101110;
DRAM[11602] = 8'b00110011;
DRAM[11603] = 8'b00101110;
DRAM[11604] = 8'b00110011;
DRAM[11605] = 8'b00110111;
DRAM[11606] = 8'b00110110;
DRAM[11607] = 8'b01000111;
DRAM[11608] = 8'b01000111;
DRAM[11609] = 8'b01010001;
DRAM[11610] = 8'b01000011;
DRAM[11611] = 8'b01010000;
DRAM[11612] = 8'b00101101;
DRAM[11613] = 8'b01001010;
DRAM[11614] = 8'b10100011;
DRAM[11615] = 8'b10010011;
DRAM[11616] = 8'b10011000;
DRAM[11617] = 8'b10010111;
DRAM[11618] = 8'b10011011;
DRAM[11619] = 8'b10011001;
DRAM[11620] = 8'b10011000;
DRAM[11621] = 8'b10011010;
DRAM[11622] = 8'b10010111;
DRAM[11623] = 8'b10010111;
DRAM[11624] = 8'b10010111;
DRAM[11625] = 8'b10010101;
DRAM[11626] = 8'b10010011;
DRAM[11627] = 8'b10010001;
DRAM[11628] = 8'b10010000;
DRAM[11629] = 8'b10001110;
DRAM[11630] = 8'b10001000;
DRAM[11631] = 8'b10000000;
DRAM[11632] = 8'b10000001;
DRAM[11633] = 8'b10111011;
DRAM[11634] = 8'b11010110;
DRAM[11635] = 8'b11010111;
DRAM[11636] = 8'b11010011;
DRAM[11637] = 8'b11010100;
DRAM[11638] = 8'b11010101;
DRAM[11639] = 8'b11011000;
DRAM[11640] = 8'b11010110;
DRAM[11641] = 8'b11010110;
DRAM[11642] = 8'b11010100;
DRAM[11643] = 8'b11010000;
DRAM[11644] = 8'b11001111;
DRAM[11645] = 8'b11001100;
DRAM[11646] = 8'b11001011;
DRAM[11647] = 8'b11001101;
DRAM[11648] = 8'b00110100;
DRAM[11649] = 8'b00110101;
DRAM[11650] = 8'b00110001;
DRAM[11651] = 8'b00110001;
DRAM[11652] = 8'b00111101;
DRAM[11653] = 8'b01011101;
DRAM[11654] = 8'b01011110;
DRAM[11655] = 8'b10000011;
DRAM[11656] = 8'b10010110;
DRAM[11657] = 8'b10100110;
DRAM[11658] = 8'b10110010;
DRAM[11659] = 8'b10110100;
DRAM[11660] = 8'b10110100;
DRAM[11661] = 8'b10110000;
DRAM[11662] = 8'b10100001;
DRAM[11663] = 8'b10000001;
DRAM[11664] = 8'b01001101;
DRAM[11665] = 8'b01000101;
DRAM[11666] = 8'b10000000;
DRAM[11667] = 8'b01100011;
DRAM[11668] = 8'b01011100;
DRAM[11669] = 8'b00110110;
DRAM[11670] = 8'b01110011;
DRAM[11671] = 8'b00110110;
DRAM[11672] = 8'b00101010;
DRAM[11673] = 8'b01010000;
DRAM[11674] = 8'b00110110;
DRAM[11675] = 8'b00111100;
DRAM[11676] = 8'b10010111;
DRAM[11677] = 8'b01101111;
DRAM[11678] = 8'b01110110;
DRAM[11679] = 8'b01111010;
DRAM[11680] = 8'b01001010;
DRAM[11681] = 8'b01010011;
DRAM[11682] = 8'b10000101;
DRAM[11683] = 8'b01110010;
DRAM[11684] = 8'b01100110;
DRAM[11685] = 8'b01110100;
DRAM[11686] = 8'b10011100;
DRAM[11687] = 8'b10101001;
DRAM[11688] = 8'b10110110;
DRAM[11689] = 8'b01000010;
DRAM[11690] = 8'b00110011;
DRAM[11691] = 8'b00110110;
DRAM[11692] = 8'b00110111;
DRAM[11693] = 8'b00111001;
DRAM[11694] = 8'b00101111;
DRAM[11695] = 8'b00110110;
DRAM[11696] = 8'b00101110;
DRAM[11697] = 8'b00110111;
DRAM[11698] = 8'b00111001;
DRAM[11699] = 8'b00111100;
DRAM[11700] = 8'b00111110;
DRAM[11701] = 8'b00110011;
DRAM[11702] = 8'b01000010;
DRAM[11703] = 8'b01001011;
DRAM[11704] = 8'b01000001;
DRAM[11705] = 8'b01001101;
DRAM[11706] = 8'b01100000;
DRAM[11707] = 8'b01100110;
DRAM[11708] = 8'b01101010;
DRAM[11709] = 8'b01110110;
DRAM[11710] = 8'b01111100;
DRAM[11711] = 8'b10000001;
DRAM[11712] = 8'b10000101;
DRAM[11713] = 8'b10001001;
DRAM[11714] = 8'b10001100;
DRAM[11715] = 8'b10001010;
DRAM[11716] = 8'b10000111;
DRAM[11717] = 8'b10000100;
DRAM[11718] = 8'b10000010;
DRAM[11719] = 8'b10000011;
DRAM[11720] = 8'b01111101;
DRAM[11721] = 8'b01111011;
DRAM[11722] = 8'b01111111;
DRAM[11723] = 8'b10001000;
DRAM[11724] = 8'b10010110;
DRAM[11725] = 8'b10001101;
DRAM[11726] = 8'b10001111;
DRAM[11727] = 8'b01000100;
DRAM[11728] = 8'b00101101;
DRAM[11729] = 8'b00101010;
DRAM[11730] = 8'b00110011;
DRAM[11731] = 8'b00110110;
DRAM[11732] = 8'b00111111;
DRAM[11733] = 8'b00110101;
DRAM[11734] = 8'b00110010;
DRAM[11735] = 8'b01010101;
DRAM[11736] = 8'b01001100;
DRAM[11737] = 8'b01010111;
DRAM[11738] = 8'b01000010;
DRAM[11739] = 8'b01001110;
DRAM[11740] = 8'b00110001;
DRAM[11741] = 8'b01001100;
DRAM[11742] = 8'b10100100;
DRAM[11743] = 8'b10010110;
DRAM[11744] = 8'b10010010;
DRAM[11745] = 8'b10011010;
DRAM[11746] = 8'b10011011;
DRAM[11747] = 8'b10011011;
DRAM[11748] = 8'b10011011;
DRAM[11749] = 8'b10011001;
DRAM[11750] = 8'b10011100;
DRAM[11751] = 8'b10011010;
DRAM[11752] = 8'b10011001;
DRAM[11753] = 8'b10010110;
DRAM[11754] = 8'b10010010;
DRAM[11755] = 8'b10010001;
DRAM[11756] = 8'b10010001;
DRAM[11757] = 8'b10001110;
DRAM[11758] = 8'b10001000;
DRAM[11759] = 8'b10000000;
DRAM[11760] = 8'b01111100;
DRAM[11761] = 8'b10111110;
DRAM[11762] = 8'b11011001;
DRAM[11763] = 8'b11011000;
DRAM[11764] = 8'b11010110;
DRAM[11765] = 8'b11010101;
DRAM[11766] = 8'b11011000;
DRAM[11767] = 8'b11011001;
DRAM[11768] = 8'b11010110;
DRAM[11769] = 8'b11010010;
DRAM[11770] = 8'b11001111;
DRAM[11771] = 8'b11001110;
DRAM[11772] = 8'b11010000;
DRAM[11773] = 8'b11010000;
DRAM[11774] = 8'b11010001;
DRAM[11775] = 8'b11010011;
DRAM[11776] = 8'b00110110;
DRAM[11777] = 8'b00110100;
DRAM[11778] = 8'b00110001;
DRAM[11779] = 8'b00101111;
DRAM[11780] = 8'b01000101;
DRAM[11781] = 8'b01100101;
DRAM[11782] = 8'b01100111;
DRAM[11783] = 8'b10000010;
DRAM[11784] = 8'b10010011;
DRAM[11785] = 8'b10100111;
DRAM[11786] = 8'b10110000;
DRAM[11787] = 8'b10110001;
DRAM[11788] = 8'b10110011;
DRAM[11789] = 8'b10110001;
DRAM[11790] = 8'b10100001;
DRAM[11791] = 8'b10000110;
DRAM[11792] = 8'b01010010;
DRAM[11793] = 8'b01000100;
DRAM[11794] = 8'b01111100;
DRAM[11795] = 8'b01100001;
DRAM[11796] = 8'b01010010;
DRAM[11797] = 8'b01000110;
DRAM[11798] = 8'b01001101;
DRAM[11799] = 8'b00110111;
DRAM[11800] = 8'b00101001;
DRAM[11801] = 8'b01010101;
DRAM[11802] = 8'b00111100;
DRAM[11803] = 8'b00110011;
DRAM[11804] = 8'b10001111;
DRAM[11805] = 8'b01111111;
DRAM[11806] = 8'b01101100;
DRAM[11807] = 8'b10000110;
DRAM[11808] = 8'b01110000;
DRAM[11809] = 8'b01011110;
DRAM[11810] = 8'b01100100;
DRAM[11811] = 8'b01101011;
DRAM[11812] = 8'b01011111;
DRAM[11813] = 8'b01101111;
DRAM[11814] = 8'b10101011;
DRAM[11815] = 8'b11001011;
DRAM[11816] = 8'b01010101;
DRAM[11817] = 8'b00110000;
DRAM[11818] = 8'b00110010;
DRAM[11819] = 8'b00110010;
DRAM[11820] = 8'b00110110;
DRAM[11821] = 8'b00111010;
DRAM[11822] = 8'b00110000;
DRAM[11823] = 8'b00110101;
DRAM[11824] = 8'b00110100;
DRAM[11825] = 8'b00110010;
DRAM[11826] = 8'b00110111;
DRAM[11827] = 8'b00110111;
DRAM[11828] = 8'b00111111;
DRAM[11829] = 8'b00110110;
DRAM[11830] = 8'b00111001;
DRAM[11831] = 8'b00111100;
DRAM[11832] = 8'b00111000;
DRAM[11833] = 8'b01000101;
DRAM[11834] = 8'b01010100;
DRAM[11835] = 8'b01011111;
DRAM[11836] = 8'b01101010;
DRAM[11837] = 8'b01110001;
DRAM[11838] = 8'b01111111;
DRAM[11839] = 8'b01111111;
DRAM[11840] = 8'b10000011;
DRAM[11841] = 8'b10001000;
DRAM[11842] = 8'b10001010;
DRAM[11843] = 8'b10001011;
DRAM[11844] = 8'b10001011;
DRAM[11845] = 8'b10001110;
DRAM[11846] = 8'b10001101;
DRAM[11847] = 8'b10010111;
DRAM[11848] = 8'b10011110;
DRAM[11849] = 8'b10100001;
DRAM[11850] = 8'b10011011;
DRAM[11851] = 8'b10011011;
DRAM[11852] = 8'b10010110;
DRAM[11853] = 8'b10010000;
DRAM[11854] = 8'b01011110;
DRAM[11855] = 8'b00111001;
DRAM[11856] = 8'b00101111;
DRAM[11857] = 8'b00101110;
DRAM[11858] = 8'b00110010;
DRAM[11859] = 8'b00110101;
DRAM[11860] = 8'b00111010;
DRAM[11861] = 8'b00110101;
DRAM[11862] = 8'b00101111;
DRAM[11863] = 8'b01010110;
DRAM[11864] = 8'b01001010;
DRAM[11865] = 8'b01010100;
DRAM[11866] = 8'b01000111;
DRAM[11867] = 8'b01001111;
DRAM[11868] = 8'b00110101;
DRAM[11869] = 8'b01000110;
DRAM[11870] = 8'b10100100;
DRAM[11871] = 8'b10011001;
DRAM[11872] = 8'b10010001;
DRAM[11873] = 8'b10011011;
DRAM[11874] = 8'b10011100;
DRAM[11875] = 8'b10011010;
DRAM[11876] = 8'b10011001;
DRAM[11877] = 8'b10011001;
DRAM[11878] = 8'b10011000;
DRAM[11879] = 8'b10010111;
DRAM[11880] = 8'b10011001;
DRAM[11881] = 8'b10010100;
DRAM[11882] = 8'b10010101;
DRAM[11883] = 8'b10010001;
DRAM[11884] = 8'b10010000;
DRAM[11885] = 8'b10001101;
DRAM[11886] = 8'b10000110;
DRAM[11887] = 8'b01111011;
DRAM[11888] = 8'b01111001;
DRAM[11889] = 8'b11000011;
DRAM[11890] = 8'b11011010;
DRAM[11891] = 8'b11011010;
DRAM[11892] = 8'b11010110;
DRAM[11893] = 8'b11010111;
DRAM[11894] = 8'b11010111;
DRAM[11895] = 8'b11010110;
DRAM[11896] = 8'b11010011;
DRAM[11897] = 8'b11010010;
DRAM[11898] = 8'b11010011;
DRAM[11899] = 8'b11010011;
DRAM[11900] = 8'b11010011;
DRAM[11901] = 8'b11010010;
DRAM[11902] = 8'b11010010;
DRAM[11903] = 8'b11010000;
DRAM[11904] = 8'b00110001;
DRAM[11905] = 8'b00110001;
DRAM[11906] = 8'b00110001;
DRAM[11907] = 8'b00110010;
DRAM[11908] = 8'b01010000;
DRAM[11909] = 8'b01101001;
DRAM[11910] = 8'b01101000;
DRAM[11911] = 8'b10000101;
DRAM[11912] = 8'b10010011;
DRAM[11913] = 8'b10100101;
DRAM[11914] = 8'b10110000;
DRAM[11915] = 8'b10101111;
DRAM[11916] = 8'b10110010;
DRAM[11917] = 8'b10110000;
DRAM[11918] = 8'b10011110;
DRAM[11919] = 8'b10000010;
DRAM[11920] = 8'b01010110;
DRAM[11921] = 8'b01000110;
DRAM[11922] = 8'b01100110;
DRAM[11923] = 8'b01100110;
DRAM[11924] = 8'b01001001;
DRAM[11925] = 8'b01010000;
DRAM[11926] = 8'b01001100;
DRAM[11927] = 8'b00110100;
DRAM[11928] = 8'b00101010;
DRAM[11929] = 8'b01010101;
DRAM[11930] = 8'b00110010;
DRAM[11931] = 8'b00111111;
DRAM[11932] = 8'b01101100;
DRAM[11933] = 8'b01100100;
DRAM[11934] = 8'b01110001;
DRAM[11935] = 8'b01111100;
DRAM[11936] = 8'b01110100;
DRAM[11937] = 8'b01100111;
DRAM[11938] = 8'b01001000;
DRAM[11939] = 8'b01111001;
DRAM[11940] = 8'b10001011;
DRAM[11941] = 8'b01010100;
DRAM[11942] = 8'b10000111;
DRAM[11943] = 8'b10000001;
DRAM[11944] = 8'b00110101;
DRAM[11945] = 8'b00101110;
DRAM[11946] = 8'b00110100;
DRAM[11947] = 8'b00110001;
DRAM[11948] = 8'b00111010;
DRAM[11949] = 8'b00111011;
DRAM[11950] = 8'b00101110;
DRAM[11951] = 8'b00111001;
DRAM[11952] = 8'b00110011;
DRAM[11953] = 8'b00110100;
DRAM[11954] = 8'b00110001;
DRAM[11955] = 8'b00110111;
DRAM[11956] = 8'b00111001;
DRAM[11957] = 8'b00110111;
DRAM[11958] = 8'b00110110;
DRAM[11959] = 8'b00111101;
DRAM[11960] = 8'b00111011;
DRAM[11961] = 8'b01000111;
DRAM[11962] = 8'b00111010;
DRAM[11963] = 8'b01001111;
DRAM[11964] = 8'b01011110;
DRAM[11965] = 8'b01101010;
DRAM[11966] = 8'b01110101;
DRAM[11967] = 8'b10000010;
DRAM[11968] = 8'b10000110;
DRAM[11969] = 8'b10001001;
DRAM[11970] = 8'b10001010;
DRAM[11971] = 8'b10001111;
DRAM[11972] = 8'b10010011;
DRAM[11973] = 8'b10011100;
DRAM[11974] = 8'b10011100;
DRAM[11975] = 8'b10100000;
DRAM[11976] = 8'b10101010;
DRAM[11977] = 8'b10101010;
DRAM[11978] = 8'b10100110;
DRAM[11979] = 8'b10011110;
DRAM[11980] = 8'b10010101;
DRAM[11981] = 8'b10010100;
DRAM[11982] = 8'b00101110;
DRAM[11983] = 8'b00111010;
DRAM[11984] = 8'b00101010;
DRAM[11985] = 8'b00101111;
DRAM[11986] = 8'b00111010;
DRAM[11987] = 8'b00111011;
DRAM[11988] = 8'b00111011;
DRAM[11989] = 8'b00110011;
DRAM[11990] = 8'b00110010;
DRAM[11991] = 8'b01011100;
DRAM[11992] = 8'b01001010;
DRAM[11993] = 8'b01100000;
DRAM[11994] = 8'b01000011;
DRAM[11995] = 8'b01001010;
DRAM[11996] = 8'b01000101;
DRAM[11997] = 8'b00111011;
DRAM[11998] = 8'b10100101;
DRAM[11999] = 8'b10011100;
DRAM[12000] = 8'b10010010;
DRAM[12001] = 8'b10011100;
DRAM[12002] = 8'b10011100;
DRAM[12003] = 8'b10011011;
DRAM[12004] = 8'b10011001;
DRAM[12005] = 8'b10010110;
DRAM[12006] = 8'b10010111;
DRAM[12007] = 8'b10010111;
DRAM[12008] = 8'b10011001;
DRAM[12009] = 8'b10010101;
DRAM[12010] = 8'b10010100;
DRAM[12011] = 8'b10010000;
DRAM[12012] = 8'b10001101;
DRAM[12013] = 8'b10001011;
DRAM[12014] = 8'b10000101;
DRAM[12015] = 8'b01111010;
DRAM[12016] = 8'b01111111;
DRAM[12017] = 8'b11001011;
DRAM[12018] = 8'b11011011;
DRAM[12019] = 8'b11011010;
DRAM[12020] = 8'b11010110;
DRAM[12021] = 8'b11010100;
DRAM[12022] = 8'b11010011;
DRAM[12023] = 8'b11010110;
DRAM[12024] = 8'b11010110;
DRAM[12025] = 8'b11010100;
DRAM[12026] = 8'b11010100;
DRAM[12027] = 8'b11010010;
DRAM[12028] = 8'b11001111;
DRAM[12029] = 8'b11001111;
DRAM[12030] = 8'b11001111;
DRAM[12031] = 8'b11001011;
DRAM[12032] = 8'b00110001;
DRAM[12033] = 8'b00110100;
DRAM[12034] = 8'b00101110;
DRAM[12035] = 8'b00110011;
DRAM[12036] = 8'b01001110;
DRAM[12037] = 8'b01100001;
DRAM[12038] = 8'b01100111;
DRAM[12039] = 8'b10000101;
DRAM[12040] = 8'b10010011;
DRAM[12041] = 8'b10100111;
DRAM[12042] = 8'b10110000;
DRAM[12043] = 8'b10110000;
DRAM[12044] = 8'b10110000;
DRAM[12045] = 8'b10101110;
DRAM[12046] = 8'b10100010;
DRAM[12047] = 8'b10000100;
DRAM[12048] = 8'b01010000;
DRAM[12049] = 8'b01000111;
DRAM[12050] = 8'b01011111;
DRAM[12051] = 8'b01011110;
DRAM[12052] = 8'b00111110;
DRAM[12053] = 8'b00111110;
DRAM[12054] = 8'b01010100;
DRAM[12055] = 8'b00111011;
DRAM[12056] = 8'b00101101;
DRAM[12057] = 8'b01001110;
DRAM[12058] = 8'b00110110;
DRAM[12059] = 8'b01000000;
DRAM[12060] = 8'b01101100;
DRAM[12061] = 8'b01010000;
DRAM[12062] = 8'b00111100;
DRAM[12063] = 8'b01101111;
DRAM[12064] = 8'b10000111;
DRAM[12065] = 8'b01111011;
DRAM[12066] = 8'b01101001;
DRAM[12067] = 8'b10000100;
DRAM[12068] = 8'b10001111;
DRAM[12069] = 8'b01010111;
DRAM[12070] = 8'b01011011;
DRAM[12071] = 8'b01100011;
DRAM[12072] = 8'b01000000;
DRAM[12073] = 8'b00110100;
DRAM[12074] = 8'b00110100;
DRAM[12075] = 8'b00110101;
DRAM[12076] = 8'b00111000;
DRAM[12077] = 8'b00111100;
DRAM[12078] = 8'b00101111;
DRAM[12079] = 8'b00111011;
DRAM[12080] = 8'b00110000;
DRAM[12081] = 8'b00110110;
DRAM[12082] = 8'b00101100;
DRAM[12083] = 8'b00110001;
DRAM[12084] = 8'b00111001;
DRAM[12085] = 8'b00110111;
DRAM[12086] = 8'b00110111;
DRAM[12087] = 8'b00111011;
DRAM[12088] = 8'b01000010;
DRAM[12089] = 8'b00111111;
DRAM[12090] = 8'b00111101;
DRAM[12091] = 8'b00110001;
DRAM[12092] = 8'b01000100;
DRAM[12093] = 8'b01010111;
DRAM[12094] = 8'b01101100;
DRAM[12095] = 8'b01111011;
DRAM[12096] = 8'b10000000;
DRAM[12097] = 8'b10000101;
DRAM[12098] = 8'b10001011;
DRAM[12099] = 8'b10010001;
DRAM[12100] = 8'b10010101;
DRAM[12101] = 8'b10011101;
DRAM[12102] = 8'b10101001;
DRAM[12103] = 8'b10100100;
DRAM[12104] = 8'b10101000;
DRAM[12105] = 8'b10100110;
DRAM[12106] = 8'b10101110;
DRAM[12107] = 8'b10100010;
DRAM[12108] = 8'b10010100;
DRAM[12109] = 8'b01111010;
DRAM[12110] = 8'b00101101;
DRAM[12111] = 8'b00111100;
DRAM[12112] = 8'b00110011;
DRAM[12113] = 8'b00110010;
DRAM[12114] = 8'b00110111;
DRAM[12115] = 8'b00111010;
DRAM[12116] = 8'b00110010;
DRAM[12117] = 8'b00110111;
DRAM[12118] = 8'b00110110;
DRAM[12119] = 8'b01100010;
DRAM[12120] = 8'b01001010;
DRAM[12121] = 8'b01100010;
DRAM[12122] = 8'b01001000;
DRAM[12123] = 8'b01000110;
DRAM[12124] = 8'b01001010;
DRAM[12125] = 8'b00111010;
DRAM[12126] = 8'b10101100;
DRAM[12127] = 8'b10100000;
DRAM[12128] = 8'b10010001;
DRAM[12129] = 8'b10011010;
DRAM[12130] = 8'b10011011;
DRAM[12131] = 8'b10010110;
DRAM[12132] = 8'b10011000;
DRAM[12133] = 8'b10010110;
DRAM[12134] = 8'b10010100;
DRAM[12135] = 8'b10010100;
DRAM[12136] = 8'b10010110;
DRAM[12137] = 8'b10010011;
DRAM[12138] = 8'b10010010;
DRAM[12139] = 8'b10001110;
DRAM[12140] = 8'b10001100;
DRAM[12141] = 8'b10001001;
DRAM[12142] = 8'b10000011;
DRAM[12143] = 8'b01111000;
DRAM[12144] = 8'b10001100;
DRAM[12145] = 8'b11010010;
DRAM[12146] = 8'b11011100;
DRAM[12147] = 8'b11011001;
DRAM[12148] = 8'b11010001;
DRAM[12149] = 8'b11010100;
DRAM[12150] = 8'b11010110;
DRAM[12151] = 8'b11010111;
DRAM[12152] = 8'b11010110;
DRAM[12153] = 8'b11010010;
DRAM[12154] = 8'b11001110;
DRAM[12155] = 8'b11001101;
DRAM[12156] = 8'b11001101;
DRAM[12157] = 8'b11001101;
DRAM[12158] = 8'b11001000;
DRAM[12159] = 8'b10111111;
DRAM[12160] = 8'b00101111;
DRAM[12161] = 8'b00110000;
DRAM[12162] = 8'b00101100;
DRAM[12163] = 8'b00101111;
DRAM[12164] = 8'b00111111;
DRAM[12165] = 8'b01011100;
DRAM[12166] = 8'b01110000;
DRAM[12167] = 8'b10000101;
DRAM[12168] = 8'b10010111;
DRAM[12169] = 8'b10100110;
DRAM[12170] = 8'b10101101;
DRAM[12171] = 8'b10110000;
DRAM[12172] = 8'b10110001;
DRAM[12173] = 8'b10110000;
DRAM[12174] = 8'b10100010;
DRAM[12175] = 8'b10000101;
DRAM[12176] = 8'b01001111;
DRAM[12177] = 8'b01000100;
DRAM[12178] = 8'b01100111;
DRAM[12179] = 8'b00111100;
DRAM[12180] = 8'b00110010;
DRAM[12181] = 8'b01001110;
DRAM[12182] = 8'b01001011;
DRAM[12183] = 8'b00111000;
DRAM[12184] = 8'b00111101;
DRAM[12185] = 8'b01000110;
DRAM[12186] = 8'b00101111;
DRAM[12187] = 8'b00110001;
DRAM[12188] = 8'b10000010;
DRAM[12189] = 8'b01100110;
DRAM[12190] = 8'b01000100;
DRAM[12191] = 8'b01010110;
DRAM[12192] = 8'b01101011;
DRAM[12193] = 8'b01111010;
DRAM[12194] = 8'b10001010;
DRAM[12195] = 8'b01111000;
DRAM[12196] = 8'b10010100;
DRAM[12197] = 8'b01100110;
DRAM[12198] = 8'b01100101;
DRAM[12199] = 8'b01000000;
DRAM[12200] = 8'b00110101;
DRAM[12201] = 8'b00110010;
DRAM[12202] = 8'b00110010;
DRAM[12203] = 8'b00110011;
DRAM[12204] = 8'b00111101;
DRAM[12205] = 8'b01000000;
DRAM[12206] = 8'b00110001;
DRAM[12207] = 8'b00111011;
DRAM[12208] = 8'b00110000;
DRAM[12209] = 8'b00110100;
DRAM[12210] = 8'b00110011;
DRAM[12211] = 8'b00110100;
DRAM[12212] = 8'b00110110;
DRAM[12213] = 8'b00111001;
DRAM[12214] = 8'b00111001;
DRAM[12215] = 8'b00111010;
DRAM[12216] = 8'b00111011;
DRAM[12217] = 8'b00111010;
DRAM[12218] = 8'b01000111;
DRAM[12219] = 8'b00110001;
DRAM[12220] = 8'b00101101;
DRAM[12221] = 8'b00111101;
DRAM[12222] = 8'b01010100;
DRAM[12223] = 8'b01100111;
DRAM[12224] = 8'b01101100;
DRAM[12225] = 8'b01111100;
DRAM[12226] = 8'b10000000;
DRAM[12227] = 8'b10001010;
DRAM[12228] = 8'b10010000;
DRAM[12229] = 8'b10010111;
DRAM[12230] = 8'b10011101;
DRAM[12231] = 8'b10101000;
DRAM[12232] = 8'b10101001;
DRAM[12233] = 8'b10100011;
DRAM[12234] = 8'b10100000;
DRAM[12235] = 8'b10011101;
DRAM[12236] = 8'b10010000;
DRAM[12237] = 8'b01101011;
DRAM[12238] = 8'b00101110;
DRAM[12239] = 8'b00111001;
DRAM[12240] = 8'b00111001;
DRAM[12241] = 8'b00110110;
DRAM[12242] = 8'b00111010;
DRAM[12243] = 8'b01000011;
DRAM[12244] = 8'b00111001;
DRAM[12245] = 8'b00110100;
DRAM[12246] = 8'b00110111;
DRAM[12247] = 8'b01100000;
DRAM[12248] = 8'b01010000;
DRAM[12249] = 8'b01011110;
DRAM[12250] = 8'b01010010;
DRAM[12251] = 8'b01001101;
DRAM[12252] = 8'b01001010;
DRAM[12253] = 8'b00111100;
DRAM[12254] = 8'b10100111;
DRAM[12255] = 8'b10011101;
DRAM[12256] = 8'b10001100;
DRAM[12257] = 8'b10010000;
DRAM[12258] = 8'b10010010;
DRAM[12259] = 8'b10010100;
DRAM[12260] = 8'b10010101;
DRAM[12261] = 8'b10010101;
DRAM[12262] = 8'b10010100;
DRAM[12263] = 8'b10010100;
DRAM[12264] = 8'b10010110;
DRAM[12265] = 8'b10010001;
DRAM[12266] = 8'b10010000;
DRAM[12267] = 8'b10001100;
DRAM[12268] = 8'b10001010;
DRAM[12269] = 8'b10001000;
DRAM[12270] = 8'b10000001;
DRAM[12271] = 8'b01110111;
DRAM[12272] = 8'b10011000;
DRAM[12273] = 8'b11010011;
DRAM[12274] = 8'b11011101;
DRAM[12275] = 8'b11010111;
DRAM[12276] = 8'b11010011;
DRAM[12277] = 8'b11010100;
DRAM[12278] = 8'b11010101;
DRAM[12279] = 8'b11010110;
DRAM[12280] = 8'b11010100;
DRAM[12281] = 8'b11001111;
DRAM[12282] = 8'b11001110;
DRAM[12283] = 8'b11001011;
DRAM[12284] = 8'b11000000;
DRAM[12285] = 8'b10101000;
DRAM[12286] = 8'b01111010;
DRAM[12287] = 8'b01001111;
DRAM[12288] = 8'b00101011;
DRAM[12289] = 8'b00110101;
DRAM[12290] = 8'b00101011;
DRAM[12291] = 8'b00101010;
DRAM[12292] = 8'b00110110;
DRAM[12293] = 8'b01011010;
DRAM[12294] = 8'b01100010;
DRAM[12295] = 8'b10000011;
DRAM[12296] = 8'b10011001;
DRAM[12297] = 8'b10100111;
DRAM[12298] = 8'b10101101;
DRAM[12299] = 8'b10101110;
DRAM[12300] = 8'b10110001;
DRAM[12301] = 8'b10110000;
DRAM[12302] = 8'b10011110;
DRAM[12303] = 8'b01111111;
DRAM[12304] = 8'b01001000;
DRAM[12305] = 8'b01110000;
DRAM[12306] = 8'b10000100;
DRAM[12307] = 8'b01110001;
DRAM[12308] = 8'b00101101;
DRAM[12309] = 8'b01001110;
DRAM[12310] = 8'b00111110;
DRAM[12311] = 8'b01000000;
DRAM[12312] = 8'b01000010;
DRAM[12313] = 8'b00110111;
DRAM[12314] = 8'b00101111;
DRAM[12315] = 8'b00110010;
DRAM[12316] = 8'b10000000;
DRAM[12317] = 8'b10000001;
DRAM[12318] = 8'b01011010;
DRAM[12319] = 8'b01000011;
DRAM[12320] = 8'b01101110;
DRAM[12321] = 8'b01101101;
DRAM[12322] = 8'b01101101;
DRAM[12323] = 8'b01111010;
DRAM[12324] = 8'b10010110;
DRAM[12325] = 8'b10000101;
DRAM[12326] = 8'b10010110;
DRAM[12327] = 8'b01111001;
DRAM[12328] = 8'b00101111;
DRAM[12329] = 8'b00110001;
DRAM[12330] = 8'b00110101;
DRAM[12331] = 8'b00110100;
DRAM[12332] = 8'b01001000;
DRAM[12333] = 8'b01000010;
DRAM[12334] = 8'b00101100;
DRAM[12335] = 8'b00111100;
DRAM[12336] = 8'b00110000;
DRAM[12337] = 8'b00110011;
DRAM[12338] = 8'b00110010;
DRAM[12339] = 8'b00110001;
DRAM[12340] = 8'b00101111;
DRAM[12341] = 8'b00111000;
DRAM[12342] = 8'b00111101;
DRAM[12343] = 8'b00111100;
DRAM[12344] = 8'b00111111;
DRAM[12345] = 8'b00110111;
DRAM[12346] = 8'b01000100;
DRAM[12347] = 8'b01001011;
DRAM[12348] = 8'b00111111;
DRAM[12349] = 8'b01000111;
DRAM[12350] = 8'b01001110;
DRAM[12351] = 8'b01010100;
DRAM[12352] = 8'b01100001;
DRAM[12353] = 8'b01101000;
DRAM[12354] = 8'b01110011;
DRAM[12355] = 8'b01111110;
DRAM[12356] = 8'b10001010;
DRAM[12357] = 8'b10010010;
DRAM[12358] = 8'b10010110;
DRAM[12359] = 8'b10011110;
DRAM[12360] = 8'b10100101;
DRAM[12361] = 8'b10011110;
DRAM[12362] = 8'b10011101;
DRAM[12363] = 8'b10001011;
DRAM[12364] = 8'b10001000;
DRAM[12365] = 8'b01010110;
DRAM[12366] = 8'b00110101;
DRAM[12367] = 8'b00110101;
DRAM[12368] = 8'b00111001;
DRAM[12369] = 8'b00111011;
DRAM[12370] = 8'b00111000;
DRAM[12371] = 8'b01000011;
DRAM[12372] = 8'b00110111;
DRAM[12373] = 8'b00110101;
DRAM[12374] = 8'b00111011;
DRAM[12375] = 8'b01100001;
DRAM[12376] = 8'b01010110;
DRAM[12377] = 8'b01011010;
DRAM[12378] = 8'b01010011;
DRAM[12379] = 8'b01010010;
DRAM[12380] = 8'b01001110;
DRAM[12381] = 8'b01001011;
DRAM[12382] = 8'b10100101;
DRAM[12383] = 8'b10010111;
DRAM[12384] = 8'b01110111;
DRAM[12385] = 8'b01110111;
DRAM[12386] = 8'b10000010;
DRAM[12387] = 8'b10000111;
DRAM[12388] = 8'b10001101;
DRAM[12389] = 8'b10001101;
DRAM[12390] = 8'b10010011;
DRAM[12391] = 8'b10010010;
DRAM[12392] = 8'b10010100;
DRAM[12393] = 8'b10001111;
DRAM[12394] = 8'b10001111;
DRAM[12395] = 8'b10001111;
DRAM[12396] = 8'b10001010;
DRAM[12397] = 8'b10000110;
DRAM[12398] = 8'b01111110;
DRAM[12399] = 8'b01110100;
DRAM[12400] = 8'b10101101;
DRAM[12401] = 8'b11011000;
DRAM[12402] = 8'b11011001;
DRAM[12403] = 8'b11010100;
DRAM[12404] = 8'b11010011;
DRAM[12405] = 8'b11010010;
DRAM[12406] = 8'b11010010;
DRAM[12407] = 8'b11010010;
DRAM[12408] = 8'b11010000;
DRAM[12409] = 8'b11001001;
DRAM[12410] = 8'b10111100;
DRAM[12411] = 8'b10100001;
DRAM[12412] = 8'b01101000;
DRAM[12413] = 8'b00110011;
DRAM[12414] = 8'b00101010;
DRAM[12415] = 8'b00101110;
DRAM[12416] = 8'b00110011;
DRAM[12417] = 8'b00110101;
DRAM[12418] = 8'b00101011;
DRAM[12419] = 8'b00101010;
DRAM[12420] = 8'b00110011;
DRAM[12421] = 8'b01001111;
DRAM[12422] = 8'b01010001;
DRAM[12423] = 8'b01111101;
DRAM[12424] = 8'b10010101;
DRAM[12425] = 8'b10100110;
DRAM[12426] = 8'b10101100;
DRAM[12427] = 8'b10101110;
DRAM[12428] = 8'b10101011;
DRAM[12429] = 8'b10101110;
DRAM[12430] = 8'b10011101;
DRAM[12431] = 8'b01111010;
DRAM[12432] = 8'b10010000;
DRAM[12433] = 8'b10010111;
DRAM[12434] = 8'b01001001;
DRAM[12435] = 8'b01101010;
DRAM[12436] = 8'b00101000;
DRAM[12437] = 8'b01001000;
DRAM[12438] = 8'b00111111;
DRAM[12439] = 8'b01000010;
DRAM[12440] = 8'b00111101;
DRAM[12441] = 8'b00111011;
DRAM[12442] = 8'b00101110;
DRAM[12443] = 8'b00101110;
DRAM[12444] = 8'b01110011;
DRAM[12445] = 8'b10000100;
DRAM[12446] = 8'b01101001;
DRAM[12447] = 8'b01000100;
DRAM[12448] = 8'b00111111;
DRAM[12449] = 8'b01011111;
DRAM[12450] = 8'b10001100;
DRAM[12451] = 8'b01100000;
DRAM[12452] = 8'b10010011;
DRAM[12453] = 8'b10000010;
DRAM[12454] = 8'b01000110;
DRAM[12455] = 8'b10010101;
DRAM[12456] = 8'b10000100;
DRAM[12457] = 8'b00101000;
DRAM[12458] = 8'b00101110;
DRAM[12459] = 8'b00110001;
DRAM[12460] = 8'b01000000;
DRAM[12461] = 8'b01000101;
DRAM[12462] = 8'b00100111;
DRAM[12463] = 8'b01000000;
DRAM[12464] = 8'b00110010;
DRAM[12465] = 8'b00110010;
DRAM[12466] = 8'b00110100;
DRAM[12467] = 8'b00110011;
DRAM[12468] = 8'b00110010;
DRAM[12469] = 8'b00110100;
DRAM[12470] = 8'b00111001;
DRAM[12471] = 8'b00110111;
DRAM[12472] = 8'b00111100;
DRAM[12473] = 8'b00110011;
DRAM[12474] = 8'b00111100;
DRAM[12475] = 8'b01001100;
DRAM[12476] = 8'b01011100;
DRAM[12477] = 8'b01101111;
DRAM[12478] = 8'b01111011;
DRAM[12479] = 8'b10000011;
DRAM[12480] = 8'b10000101;
DRAM[12481] = 8'b10001011;
DRAM[12482] = 8'b10001000;
DRAM[12483] = 8'b10001110;
DRAM[12484] = 8'b10001111;
DRAM[12485] = 8'b10011000;
DRAM[12486] = 8'b10011100;
DRAM[12487] = 8'b10011011;
DRAM[12488] = 8'b10011110;
DRAM[12489] = 8'b10011111;
DRAM[12490] = 8'b10100011;
DRAM[12491] = 8'b10101110;
DRAM[12492] = 8'b10111100;
DRAM[12493] = 8'b10110011;
DRAM[12494] = 8'b10001000;
DRAM[12495] = 8'b01001100;
DRAM[12496] = 8'b00110100;
DRAM[12497] = 8'b00110101;
DRAM[12498] = 8'b00110100;
DRAM[12499] = 8'b00111000;
DRAM[12500] = 8'b00110010;
DRAM[12501] = 8'b00110110;
DRAM[12502] = 8'b00111010;
DRAM[12503] = 8'b01011101;
DRAM[12504] = 8'b01010010;
DRAM[12505] = 8'b01011110;
DRAM[12506] = 8'b01001111;
DRAM[12507] = 8'b01010010;
DRAM[12508] = 8'b01000111;
DRAM[12509] = 8'b01010100;
DRAM[12510] = 8'b10100010;
DRAM[12511] = 8'b10001101;
DRAM[12512] = 8'b01101111;
DRAM[12513] = 8'b01101111;
DRAM[12514] = 8'b01110001;
DRAM[12515] = 8'b01110101;
DRAM[12516] = 8'b01111000;
DRAM[12517] = 8'b01111011;
DRAM[12518] = 8'b01111110;
DRAM[12519] = 8'b10000010;
DRAM[12520] = 8'b10001011;
DRAM[12521] = 8'b10001111;
DRAM[12522] = 8'b10001101;
DRAM[12523] = 8'b10001011;
DRAM[12524] = 8'b10001001;
DRAM[12525] = 8'b10000001;
DRAM[12526] = 8'b01111100;
DRAM[12527] = 8'b01110100;
DRAM[12528] = 8'b11000000;
DRAM[12529] = 8'b11011000;
DRAM[12530] = 8'b11010100;
DRAM[12531] = 8'b11010001;
DRAM[12532] = 8'b11010000;
DRAM[12533] = 8'b11010001;
DRAM[12534] = 8'b11010000;
DRAM[12535] = 8'b11001101;
DRAM[12536] = 8'b11001000;
DRAM[12537] = 8'b10110010;
DRAM[12538] = 8'b10001100;
DRAM[12539] = 8'b01000000;
DRAM[12540] = 8'b00101000;
DRAM[12541] = 8'b00101011;
DRAM[12542] = 8'b00110111;
DRAM[12543] = 8'b01000100;
DRAM[12544] = 8'b01000010;
DRAM[12545] = 8'b00111101;
DRAM[12546] = 8'b00110011;
DRAM[12547] = 8'b00101111;
DRAM[12548] = 8'b00110001;
DRAM[12549] = 8'b01000110;
DRAM[12550] = 8'b01001010;
DRAM[12551] = 8'b01110110;
DRAM[12552] = 8'b10010000;
DRAM[12553] = 8'b10100100;
DRAM[12554] = 8'b10101010;
DRAM[12555] = 8'b10101011;
DRAM[12556] = 8'b10101100;
DRAM[12557] = 8'b10101110;
DRAM[12558] = 8'b10011011;
DRAM[12559] = 8'b10100110;
DRAM[12560] = 8'b01111000;
DRAM[12561] = 8'b01001001;
DRAM[12562] = 8'b01000110;
DRAM[12563] = 8'b01011000;
DRAM[12564] = 8'b00101010;
DRAM[12565] = 8'b01000000;
DRAM[12566] = 8'b01001010;
DRAM[12567] = 8'b00111100;
DRAM[12568] = 8'b00110101;
DRAM[12569] = 8'b01010101;
DRAM[12570] = 8'b00111110;
DRAM[12571] = 8'b00110011;
DRAM[12572] = 8'b01010111;
DRAM[12573] = 8'b01111101;
DRAM[12574] = 8'b10000000;
DRAM[12575] = 8'b01011001;
DRAM[12576] = 8'b01000110;
DRAM[12577] = 8'b01111110;
DRAM[12578] = 8'b10000110;
DRAM[12579] = 8'b01011000;
DRAM[12580] = 8'b01100011;
DRAM[12581] = 8'b01111010;
DRAM[12582] = 8'b01011010;
DRAM[12583] = 8'b01100011;
DRAM[12584] = 8'b10010101;
DRAM[12585] = 8'b10000011;
DRAM[12586] = 8'b00101100;
DRAM[12587] = 8'b00110111;
DRAM[12588] = 8'b01001000;
DRAM[12589] = 8'b01000010;
DRAM[12590] = 8'b00101100;
DRAM[12591] = 8'b01000000;
DRAM[12592] = 8'b00110100;
DRAM[12593] = 8'b00110011;
DRAM[12594] = 8'b00110010;
DRAM[12595] = 8'b00110011;
DRAM[12596] = 8'b00110001;
DRAM[12597] = 8'b00110100;
DRAM[12598] = 8'b00110110;
DRAM[12599] = 8'b00111101;
DRAM[12600] = 8'b00111010;
DRAM[12601] = 8'b00111000;
DRAM[12602] = 8'b00110111;
DRAM[12603] = 8'b01010010;
DRAM[12604] = 8'b01101000;
DRAM[12605] = 8'b01111000;
DRAM[12606] = 8'b10000001;
DRAM[12607] = 8'b01111110;
DRAM[12608] = 8'b10000001;
DRAM[12609] = 8'b10000100;
DRAM[12610] = 8'b10000101;
DRAM[12611] = 8'b10001010;
DRAM[12612] = 8'b10001101;
DRAM[12613] = 8'b10010011;
DRAM[12614] = 8'b10010010;
DRAM[12615] = 8'b10010010;
DRAM[12616] = 8'b10010001;
DRAM[12617] = 8'b10010100;
DRAM[12618] = 8'b10100001;
DRAM[12619] = 8'b10101111;
DRAM[12620] = 8'b10111110;
DRAM[12621] = 8'b11000110;
DRAM[12622] = 8'b11001001;
DRAM[12623] = 8'b11001100;
DRAM[12624] = 8'b10011100;
DRAM[12625] = 8'b01011001;
DRAM[12626] = 8'b00110101;
DRAM[12627] = 8'b00110110;
DRAM[12628] = 8'b00101111;
DRAM[12629] = 8'b00101110;
DRAM[12630] = 8'b01000010;
DRAM[12631] = 8'b01011101;
DRAM[12632] = 8'b01010100;
DRAM[12633] = 8'b01011011;
DRAM[12634] = 8'b01001101;
DRAM[12635] = 8'b01010100;
DRAM[12636] = 8'b01001100;
DRAM[12637] = 8'b01011000;
DRAM[12638] = 8'b10100010;
DRAM[12639] = 8'b10000001;
DRAM[12640] = 8'b01111001;
DRAM[12641] = 8'b10000000;
DRAM[12642] = 8'b01110100;
DRAM[12643] = 8'b01110010;
DRAM[12644] = 8'b01110001;
DRAM[12645] = 8'b01101101;
DRAM[12646] = 8'b01101100;
DRAM[12647] = 8'b01110000;
DRAM[12648] = 8'b01110010;
DRAM[12649] = 8'b01111000;
DRAM[12650] = 8'b01111010;
DRAM[12651] = 8'b01111101;
DRAM[12652] = 8'b01111110;
DRAM[12653] = 8'b01111111;
DRAM[12654] = 8'b01110111;
DRAM[12655] = 8'b01111001;
DRAM[12656] = 8'b11000101;
DRAM[12657] = 8'b11010100;
DRAM[12658] = 8'b11001110;
DRAM[12659] = 8'b11001110;
DRAM[12660] = 8'b11010001;
DRAM[12661] = 8'b11010001;
DRAM[12662] = 8'b11010000;
DRAM[12663] = 8'b11000110;
DRAM[12664] = 8'b10111010;
DRAM[12665] = 8'b10011110;
DRAM[12666] = 8'b01010010;
DRAM[12667] = 8'b00101101;
DRAM[12668] = 8'b00110001;
DRAM[12669] = 8'b01000001;
DRAM[12670] = 8'b01010011;
DRAM[12671] = 8'b01001110;
DRAM[12672] = 8'b01110101;
DRAM[12673] = 8'b01011000;
DRAM[12674] = 8'b01000100;
DRAM[12675] = 8'b00110110;
DRAM[12676] = 8'b00111101;
DRAM[12677] = 8'b00111100;
DRAM[12678] = 8'b00111001;
DRAM[12679] = 8'b01011111;
DRAM[12680] = 8'b10001010;
DRAM[12681] = 8'b10100101;
DRAM[12682] = 8'b10101010;
DRAM[12683] = 8'b10101100;
DRAM[12684] = 8'b10101010;
DRAM[12685] = 8'b10110010;
DRAM[12686] = 8'b10101110;
DRAM[12687] = 8'b10001111;
DRAM[12688] = 8'b01001110;
DRAM[12689] = 8'b01001110;
DRAM[12690] = 8'b10000011;
DRAM[12691] = 8'b00100101;
DRAM[12692] = 8'b00100110;
DRAM[12693] = 8'b00101010;
DRAM[12694] = 8'b01001110;
DRAM[12695] = 8'b01000011;
DRAM[12696] = 8'b00101010;
DRAM[12697] = 8'b01001010;
DRAM[12698] = 8'b01010111;
DRAM[12699] = 8'b01000000;
DRAM[12700] = 8'b00111001;
DRAM[12701] = 8'b01100100;
DRAM[12702] = 8'b01110001;
DRAM[12703] = 8'b01011110;
DRAM[12704] = 8'b01101001;
DRAM[12705] = 8'b10011010;
DRAM[12706] = 8'b01010001;
DRAM[12707] = 8'b01011100;
DRAM[12708] = 8'b01101110;
DRAM[12709] = 8'b01101101;
DRAM[12710] = 8'b01100010;
DRAM[12711] = 8'b10011001;
DRAM[12712] = 8'b01110101;
DRAM[12713] = 8'b01011001;
DRAM[12714] = 8'b01010111;
DRAM[12715] = 8'b00110100;
DRAM[12716] = 8'b00111111;
DRAM[12717] = 8'b00111100;
DRAM[12718] = 8'b00101101;
DRAM[12719] = 8'b01001001;
DRAM[12720] = 8'b00110100;
DRAM[12721] = 8'b00101110;
DRAM[12722] = 8'b00110010;
DRAM[12723] = 8'b00110111;
DRAM[12724] = 8'b00110010;
DRAM[12725] = 8'b00110010;
DRAM[12726] = 8'b00110011;
DRAM[12727] = 8'b00111101;
DRAM[12728] = 8'b00111110;
DRAM[12729] = 8'b00111011;
DRAM[12730] = 8'b00110000;
DRAM[12731] = 8'b01010000;
DRAM[12732] = 8'b01101000;
DRAM[12733] = 8'b01111000;
DRAM[12734] = 8'b01111100;
DRAM[12735] = 8'b01111101;
DRAM[12736] = 8'b01111101;
DRAM[12737] = 8'b10000100;
DRAM[12738] = 8'b10000110;
DRAM[12739] = 8'b10001000;
DRAM[12740] = 8'b10001011;
DRAM[12741] = 8'b10001110;
DRAM[12742] = 8'b10001110;
DRAM[12743] = 8'b10001011;
DRAM[12744] = 8'b10001111;
DRAM[12745] = 8'b10010101;
DRAM[12746] = 8'b10100110;
DRAM[12747] = 8'b10110001;
DRAM[12748] = 8'b10111111;
DRAM[12749] = 8'b11000101;
DRAM[12750] = 8'b11001000;
DRAM[12751] = 8'b11001001;
DRAM[12752] = 8'b11001010;
DRAM[12753] = 8'b11001111;
DRAM[12754] = 8'b10101001;
DRAM[12755] = 8'b01001010;
DRAM[12756] = 8'b00101000;
DRAM[12757] = 8'b00100100;
DRAM[12758] = 8'b00111011;
DRAM[12759] = 8'b01010011;
DRAM[12760] = 8'b01010011;
DRAM[12761] = 8'b01011000;
DRAM[12762] = 8'b01000111;
DRAM[12763] = 8'b01010010;
DRAM[12764] = 8'b01000100;
DRAM[12765] = 8'b01100000;
DRAM[12766] = 8'b10010111;
DRAM[12767] = 8'b10000110;
DRAM[12768] = 8'b10000111;
DRAM[12769] = 8'b10001001;
DRAM[12770] = 8'b10000100;
DRAM[12771] = 8'b01111110;
DRAM[12772] = 8'b01111100;
DRAM[12773] = 8'b01110100;
DRAM[12774] = 8'b01101100;
DRAM[12775] = 8'b01100111;
DRAM[12776] = 8'b01100001;
DRAM[12777] = 8'b01100110;
DRAM[12778] = 8'b01100110;
DRAM[12779] = 8'b01100011;
DRAM[12780] = 8'b01101000;
DRAM[12781] = 8'b01101110;
DRAM[12782] = 8'b01100101;
DRAM[12783] = 8'b01101100;
DRAM[12784] = 8'b10111111;
DRAM[12785] = 8'b11010001;
DRAM[12786] = 8'b11001100;
DRAM[12787] = 8'b11001111;
DRAM[12788] = 8'b11010001;
DRAM[12789] = 8'b11010000;
DRAM[12790] = 8'b11001110;
DRAM[12791] = 8'b10111110;
DRAM[12792] = 8'b10001110;
DRAM[12793] = 8'b01000000;
DRAM[12794] = 8'b00110010;
DRAM[12795] = 8'b00111000;
DRAM[12796] = 8'b01000000;
DRAM[12797] = 8'b01001111;
DRAM[12798] = 8'b01010101;
DRAM[12799] = 8'b01010110;
DRAM[12800] = 8'b10000101;
DRAM[12801] = 8'b10000000;
DRAM[12802] = 8'b01100110;
DRAM[12803] = 8'b01001111;
DRAM[12804] = 8'b01001010;
DRAM[12805] = 8'b00111101;
DRAM[12806] = 8'b00110110;
DRAM[12807] = 8'b01011000;
DRAM[12808] = 8'b10000111;
DRAM[12809] = 8'b10100010;
DRAM[12810] = 8'b10101001;
DRAM[12811] = 8'b10101100;
DRAM[12812] = 8'b10101011;
DRAM[12813] = 8'b10101111;
DRAM[12814] = 8'b10100001;
DRAM[12815] = 8'b10000100;
DRAM[12816] = 8'b01011000;
DRAM[12817] = 8'b10010001;
DRAM[12818] = 8'b01011000;
DRAM[12819] = 8'b00101000;
DRAM[12820] = 8'b00101000;
DRAM[12821] = 8'b00101001;
DRAM[12822] = 8'b00111111;
DRAM[12823] = 8'b01100000;
DRAM[12824] = 8'b00100001;
DRAM[12825] = 8'b00110101;
DRAM[12826] = 8'b01100101;
DRAM[12827] = 8'b01011101;
DRAM[12828] = 8'b00110001;
DRAM[12829] = 8'b00101100;
DRAM[12830] = 8'b01101001;
DRAM[12831] = 8'b01111000;
DRAM[12832] = 8'b01100100;
DRAM[12833] = 8'b01101110;
DRAM[12834] = 8'b01001110;
DRAM[12835] = 8'b01101111;
DRAM[12836] = 8'b01101000;
DRAM[12837] = 8'b01111011;
DRAM[12838] = 8'b01110111;
DRAM[12839] = 8'b01111111;
DRAM[12840] = 8'b01111111;
DRAM[12841] = 8'b00111000;
DRAM[12842] = 8'b10001100;
DRAM[12843] = 8'b00110110;
DRAM[12844] = 8'b01000000;
DRAM[12845] = 8'b00110011;
DRAM[12846] = 8'b00101010;
DRAM[12847] = 8'b01001001;
DRAM[12848] = 8'b00110010;
DRAM[12849] = 8'b00110010;
DRAM[12850] = 8'b00101100;
DRAM[12851] = 8'b00111001;
DRAM[12852] = 8'b00111010;
DRAM[12853] = 8'b00110000;
DRAM[12854] = 8'b00110101;
DRAM[12855] = 8'b00111000;
DRAM[12856] = 8'b01000010;
DRAM[12857] = 8'b00111101;
DRAM[12858] = 8'b00110011;
DRAM[12859] = 8'b01000110;
DRAM[12860] = 8'b01100100;
DRAM[12861] = 8'b01110100;
DRAM[12862] = 8'b01111001;
DRAM[12863] = 8'b01111100;
DRAM[12864] = 8'b10000000;
DRAM[12865] = 8'b01111111;
DRAM[12866] = 8'b10000111;
DRAM[12867] = 8'b10001011;
DRAM[12868] = 8'b10001100;
DRAM[12869] = 8'b10001100;
DRAM[12870] = 8'b10001010;
DRAM[12871] = 8'b10010000;
DRAM[12872] = 8'b10010011;
DRAM[12873] = 8'b10011100;
DRAM[12874] = 8'b10100111;
DRAM[12875] = 8'b10110100;
DRAM[12876] = 8'b10111101;
DRAM[12877] = 8'b10111111;
DRAM[12878] = 8'b11000010;
DRAM[12879] = 8'b11000100;
DRAM[12880] = 8'b11001010;
DRAM[12881] = 8'b11001011;
DRAM[12882] = 8'b11010000;
DRAM[12883] = 8'b11010010;
DRAM[12884] = 8'b01111100;
DRAM[12885] = 8'b00100110;
DRAM[12886] = 8'b00111100;
DRAM[12887] = 8'b01001010;
DRAM[12888] = 8'b01010011;
DRAM[12889] = 8'b01001111;
DRAM[12890] = 8'b01000100;
DRAM[12891] = 8'b01001101;
DRAM[12892] = 8'b01000100;
DRAM[12893] = 8'b01100110;
DRAM[12894] = 8'b10010100;
DRAM[12895] = 8'b10001110;
DRAM[12896] = 8'b10001111;
DRAM[12897] = 8'b10001011;
DRAM[12898] = 8'b10001100;
DRAM[12899] = 8'b10000101;
DRAM[12900] = 8'b10000110;
DRAM[12901] = 8'b10000100;
DRAM[12902] = 8'b01111101;
DRAM[12903] = 8'b01110101;
DRAM[12904] = 8'b01101111;
DRAM[12905] = 8'b01100100;
DRAM[12906] = 8'b01011111;
DRAM[12907] = 8'b01011000;
DRAM[12908] = 8'b01100110;
DRAM[12909] = 8'b01110110;
DRAM[12910] = 8'b01100000;
DRAM[12911] = 8'b01010101;
DRAM[12912] = 8'b10111110;
DRAM[12913] = 8'b11001111;
DRAM[12914] = 8'b11001110;
DRAM[12915] = 8'b11010010;
DRAM[12916] = 8'b11010000;
DRAM[12917] = 8'b11001101;
DRAM[12918] = 8'b10111100;
DRAM[12919] = 8'b10010000;
DRAM[12920] = 8'b01000010;
DRAM[12921] = 8'b00110100;
DRAM[12922] = 8'b01001101;
DRAM[12923] = 8'b01001011;
DRAM[12924] = 8'b01010000;
DRAM[12925] = 8'b01010101;
DRAM[12926] = 8'b01011000;
DRAM[12927] = 8'b01010110;
DRAM[12928] = 8'b10000110;
DRAM[12929] = 8'b10001101;
DRAM[12930] = 8'b10000111;
DRAM[12931] = 8'b01110010;
DRAM[12932] = 8'b01011111;
DRAM[12933] = 8'b01000101;
DRAM[12934] = 8'b00110000;
DRAM[12935] = 8'b01010101;
DRAM[12936] = 8'b10000111;
DRAM[12937] = 8'b10100011;
DRAM[12938] = 8'b10101010;
DRAM[12939] = 8'b10101010;
DRAM[12940] = 8'b10101100;
DRAM[12941] = 8'b10101100;
DRAM[12942] = 8'b10011111;
DRAM[12943] = 8'b10000010;
DRAM[12944] = 8'b10110011;
DRAM[12945] = 8'b01110110;
DRAM[12946] = 8'b00101001;
DRAM[12947] = 8'b00101010;
DRAM[12948] = 8'b00101000;
DRAM[12949] = 8'b00100101;
DRAM[12950] = 8'b01100000;
DRAM[12951] = 8'b01111000;
DRAM[12952] = 8'b01010010;
DRAM[12953] = 8'b01110000;
DRAM[12954] = 8'b01010100;
DRAM[12955] = 8'b01001100;
DRAM[12956] = 8'b00110101;
DRAM[12957] = 8'b01100011;
DRAM[12958] = 8'b01000111;
DRAM[12959] = 8'b01011100;
DRAM[12960] = 8'b01101010;
DRAM[12961] = 8'b00111100;
DRAM[12962] = 8'b01001100;
DRAM[12963] = 8'b01011010;
DRAM[12964] = 8'b01111000;
DRAM[12965] = 8'b10000000;
DRAM[12966] = 8'b10001100;
DRAM[12967] = 8'b01111111;
DRAM[12968] = 8'b01001110;
DRAM[12969] = 8'b01101010;
DRAM[12970] = 8'b01000110;
DRAM[12971] = 8'b01110010;
DRAM[12972] = 8'b00110111;
DRAM[12973] = 8'b00110010;
DRAM[12974] = 8'b00101111;
DRAM[12975] = 8'b01010000;
DRAM[12976] = 8'b00111000;
DRAM[12977] = 8'b00110001;
DRAM[12978] = 8'b00110000;
DRAM[12979] = 8'b00110100;
DRAM[12980] = 8'b01000000;
DRAM[12981] = 8'b00110101;
DRAM[12982] = 8'b00110101;
DRAM[12983] = 8'b01000001;
DRAM[12984] = 8'b01000100;
DRAM[12985] = 8'b01000011;
DRAM[12986] = 8'b00110101;
DRAM[12987] = 8'b01000101;
DRAM[12988] = 8'b01100100;
DRAM[12989] = 8'b01110101;
DRAM[12990] = 8'b01111001;
DRAM[12991] = 8'b10000001;
DRAM[12992] = 8'b01111100;
DRAM[12993] = 8'b10000000;
DRAM[12994] = 8'b10001010;
DRAM[12995] = 8'b10001111;
DRAM[12996] = 8'b10001011;
DRAM[12997] = 8'b10001010;
DRAM[12998] = 8'b10001000;
DRAM[12999] = 8'b10010001;
DRAM[13000] = 8'b10010110;
DRAM[13001] = 8'b10011111;
DRAM[13002] = 8'b10101010;
DRAM[13003] = 8'b10110100;
DRAM[13004] = 8'b10111011;
DRAM[13005] = 8'b10111100;
DRAM[13006] = 8'b11000000;
DRAM[13007] = 8'b11000000;
DRAM[13008] = 8'b11000111;
DRAM[13009] = 8'b11001011;
DRAM[13010] = 8'b11001101;
DRAM[13011] = 8'b11010001;
DRAM[13012] = 8'b11010100;
DRAM[13013] = 8'b10100011;
DRAM[13014] = 8'b00110110;
DRAM[13015] = 8'b00111111;
DRAM[13016] = 8'b01001011;
DRAM[13017] = 8'b01000110;
DRAM[13018] = 8'b01000010;
DRAM[13019] = 8'b01001011;
DRAM[13020] = 8'b00111101;
DRAM[13021] = 8'b01101100;
DRAM[13022] = 8'b10010001;
DRAM[13023] = 8'b10010011;
DRAM[13024] = 8'b10010110;
DRAM[13025] = 8'b10010001;
DRAM[13026] = 8'b10010001;
DRAM[13027] = 8'b10001100;
DRAM[13028] = 8'b10001011;
DRAM[13029] = 8'b10000111;
DRAM[13030] = 8'b10000011;
DRAM[13031] = 8'b01111110;
DRAM[13032] = 8'b01111011;
DRAM[13033] = 8'b01110101;
DRAM[13034] = 8'b01101101;
DRAM[13035] = 8'b01100101;
DRAM[13036] = 8'b01110010;
DRAM[13037] = 8'b10000001;
DRAM[13038] = 8'b01100011;
DRAM[13039] = 8'b01100110;
DRAM[13040] = 8'b11000101;
DRAM[13041] = 8'b11010010;
DRAM[13042] = 8'b11010001;
DRAM[13043] = 8'b11010100;
DRAM[13044] = 8'b11010001;
DRAM[13045] = 8'b11001010;
DRAM[13046] = 8'b10000111;
DRAM[13047] = 8'b00111001;
DRAM[13048] = 8'b00110111;
DRAM[13049] = 8'b01010101;
DRAM[13050] = 8'b01001111;
DRAM[13051] = 8'b01001110;
DRAM[13052] = 8'b01011011;
DRAM[13053] = 8'b01100000;
DRAM[13054] = 8'b01011001;
DRAM[13055] = 8'b01010110;
DRAM[13056] = 8'b10000011;
DRAM[13057] = 8'b10010001;
DRAM[13058] = 8'b10010100;
DRAM[13059] = 8'b10001011;
DRAM[13060] = 8'b01110101;
DRAM[13061] = 8'b01001110;
DRAM[13062] = 8'b00101110;
DRAM[13063] = 8'b01011000;
DRAM[13064] = 8'b10001000;
DRAM[13065] = 8'b10100101;
DRAM[13066] = 8'b10101110;
DRAM[13067] = 8'b10101110;
DRAM[13068] = 8'b10101101;
DRAM[13069] = 8'b10110000;
DRAM[13070] = 8'b10011101;
DRAM[13071] = 8'b10101001;
DRAM[13072] = 8'b10100011;
DRAM[13073] = 8'b01101000;
DRAM[13074] = 8'b00111100;
DRAM[13075] = 8'b00101110;
DRAM[13076] = 8'b00110000;
DRAM[13077] = 8'b00110011;
DRAM[13078] = 8'b01000010;
DRAM[13079] = 8'b00101000;
DRAM[13080] = 8'b01001110;
DRAM[13081] = 8'b01000001;
DRAM[13082] = 8'b00111100;
DRAM[13083] = 8'b00111101;
DRAM[13084] = 8'b01010010;
DRAM[13085] = 8'b01010000;
DRAM[13086] = 8'b00101110;
DRAM[13087] = 8'b01111100;
DRAM[13088] = 8'b00111001;
DRAM[13089] = 8'b01000010;
DRAM[13090] = 8'b01000110;
DRAM[13091] = 8'b01100100;
DRAM[13092] = 8'b01100001;
DRAM[13093] = 8'b10000010;
DRAM[13094] = 8'b10000111;
DRAM[13095] = 8'b10010111;
DRAM[13096] = 8'b01000001;
DRAM[13097] = 8'b01111101;
DRAM[13098] = 8'b01011000;
DRAM[13099] = 8'b10001000;
DRAM[13100] = 8'b00110011;
DRAM[13101] = 8'b00101110;
DRAM[13102] = 8'b00101100;
DRAM[13103] = 8'b01001101;
DRAM[13104] = 8'b00110101;
DRAM[13105] = 8'b00110100;
DRAM[13106] = 8'b00110100;
DRAM[13107] = 8'b00111001;
DRAM[13108] = 8'b01000100;
DRAM[13109] = 8'b00110011;
DRAM[13110] = 8'b00110111;
DRAM[13111] = 8'b01001001;
DRAM[13112] = 8'b01000110;
DRAM[13113] = 8'b01011100;
DRAM[13114] = 8'b00110000;
DRAM[13115] = 8'b00111111;
DRAM[13116] = 8'b01100100;
DRAM[13117] = 8'b01110101;
DRAM[13118] = 8'b01111111;
DRAM[13119] = 8'b01110100;
DRAM[13120] = 8'b01111110;
DRAM[13121] = 8'b10001011;
DRAM[13122] = 8'b10001000;
DRAM[13123] = 8'b10001100;
DRAM[13124] = 8'b10001101;
DRAM[13125] = 8'b10001011;
DRAM[13126] = 8'b10001101;
DRAM[13127] = 8'b10010011;
DRAM[13128] = 8'b10011101;
DRAM[13129] = 8'b10100001;
DRAM[13130] = 8'b10100110;
DRAM[13131] = 8'b10101111;
DRAM[13132] = 8'b10110010;
DRAM[13133] = 8'b10111000;
DRAM[13134] = 8'b10111011;
DRAM[13135] = 8'b10111111;
DRAM[13136] = 8'b11000100;
DRAM[13137] = 8'b11000111;
DRAM[13138] = 8'b11001101;
DRAM[13139] = 8'b11010000;
DRAM[13140] = 8'b11010100;
DRAM[13141] = 8'b11010101;
DRAM[13142] = 8'b10101011;
DRAM[13143] = 8'b00110110;
DRAM[13144] = 8'b01000010;
DRAM[13145] = 8'b00110110;
DRAM[13146] = 8'b01001000;
DRAM[13147] = 8'b01000101;
DRAM[13148] = 8'b00111011;
DRAM[13149] = 8'b01111010;
DRAM[13150] = 8'b10001111;
DRAM[13151] = 8'b10010001;
DRAM[13152] = 8'b10010100;
DRAM[13153] = 8'b10001111;
DRAM[13154] = 8'b10010000;
DRAM[13155] = 8'b10001111;
DRAM[13156] = 8'b10001111;
DRAM[13157] = 8'b10001010;
DRAM[13158] = 8'b10001001;
DRAM[13159] = 8'b10000111;
DRAM[13160] = 8'b10000000;
DRAM[13161] = 8'b01111110;
DRAM[13162] = 8'b01111010;
DRAM[13163] = 8'b01110001;
DRAM[13164] = 8'b01111010;
DRAM[13165] = 8'b10000010;
DRAM[13166] = 8'b01101011;
DRAM[13167] = 8'b10001100;
DRAM[13168] = 8'b11001101;
DRAM[13169] = 8'b11010011;
DRAM[13170] = 8'b11010101;
DRAM[13171] = 8'b11010100;
DRAM[13172] = 8'b11001011;
DRAM[13173] = 8'b10110110;
DRAM[13174] = 8'b01011010;
DRAM[13175] = 8'b00110000;
DRAM[13176] = 8'b01010100;
DRAM[13177] = 8'b01011011;
DRAM[13178] = 8'b01010101;
DRAM[13179] = 8'b01011000;
DRAM[13180] = 8'b01100110;
DRAM[13181] = 8'b01100000;
DRAM[13182] = 8'b01011000;
DRAM[13183] = 8'b01011100;
DRAM[13184] = 8'b01101110;
DRAM[13185] = 8'b10000111;
DRAM[13186] = 8'b10010110;
DRAM[13187] = 8'b10010111;
DRAM[13188] = 8'b10010000;
DRAM[13189] = 8'b01100010;
DRAM[13190] = 8'b00110000;
DRAM[13191] = 8'b01010110;
DRAM[13192] = 8'b10001010;
DRAM[13193] = 8'b10100101;
DRAM[13194] = 8'b10110000;
DRAM[13195] = 8'b10101111;
DRAM[13196] = 8'b10110000;
DRAM[13197] = 8'b10110000;
DRAM[13198] = 8'b10011111;
DRAM[13199] = 8'b10100011;
DRAM[13200] = 8'b10010110;
DRAM[13201] = 8'b01100000;
DRAM[13202] = 8'b00100100;
DRAM[13203] = 8'b00101101;
DRAM[13204] = 8'b00110100;
DRAM[13205] = 8'b00110101;
DRAM[13206] = 8'b01000011;
DRAM[13207] = 8'b00110110;
DRAM[13208] = 8'b00111101;
DRAM[13209] = 8'b00110011;
DRAM[13210] = 8'b01001110;
DRAM[13211] = 8'b00111010;
DRAM[13212] = 8'b00101010;
DRAM[13213] = 8'b01000000;
DRAM[13214] = 8'b00101110;
DRAM[13215] = 8'b01100000;
DRAM[13216] = 8'b00111101;
DRAM[13217] = 8'b01000000;
DRAM[13218] = 8'b01001101;
DRAM[13219] = 8'b01011000;
DRAM[13220] = 8'b01100001;
DRAM[13221] = 8'b01110001;
DRAM[13222] = 8'b10001001;
DRAM[13223] = 8'b01110110;
DRAM[13224] = 8'b10000101;
DRAM[13225] = 8'b01101110;
DRAM[13226] = 8'b10000111;
DRAM[13227] = 8'b00101110;
DRAM[13228] = 8'b01110000;
DRAM[13229] = 8'b00101010;
DRAM[13230] = 8'b00101111;
DRAM[13231] = 8'b01010001;
DRAM[13232] = 8'b01000000;
DRAM[13233] = 8'b00111000;
DRAM[13234] = 8'b00110011;
DRAM[13235] = 8'b00111011;
DRAM[13236] = 8'b01000000;
DRAM[13237] = 8'b00110111;
DRAM[13238] = 8'b00111000;
DRAM[13239] = 8'b01001010;
DRAM[13240] = 8'b01001101;
DRAM[13241] = 8'b01101010;
DRAM[13242] = 8'b00111010;
DRAM[13243] = 8'b00111111;
DRAM[13244] = 8'b01101010;
DRAM[13245] = 8'b01111011;
DRAM[13246] = 8'b01110100;
DRAM[13247] = 8'b01111111;
DRAM[13248] = 8'b10000111;
DRAM[13249] = 8'b10001011;
DRAM[13250] = 8'b10001011;
DRAM[13251] = 8'b10001100;
DRAM[13252] = 8'b10001011;
DRAM[13253] = 8'b10001011;
DRAM[13254] = 8'b10001101;
DRAM[13255] = 8'b10010111;
DRAM[13256] = 8'b10011100;
DRAM[13257] = 8'b10100000;
DRAM[13258] = 8'b10100101;
DRAM[13259] = 8'b10101001;
DRAM[13260] = 8'b10101110;
DRAM[13261] = 8'b10110010;
DRAM[13262] = 8'b10110111;
DRAM[13263] = 8'b10111000;
DRAM[13264] = 8'b11000000;
DRAM[13265] = 8'b11000101;
DRAM[13266] = 8'b11001001;
DRAM[13267] = 8'b11001111;
DRAM[13268] = 8'b11010001;
DRAM[13269] = 8'b11010101;
DRAM[13270] = 8'b11011001;
DRAM[13271] = 8'b10010110;
DRAM[13272] = 8'b00110011;
DRAM[13273] = 8'b00101101;
DRAM[13274] = 8'b01000100;
DRAM[13275] = 8'b01000000;
DRAM[13276] = 8'b00110011;
DRAM[13277] = 8'b10001001;
DRAM[13278] = 8'b10001010;
DRAM[13279] = 8'b10010001;
DRAM[13280] = 8'b10010110;
DRAM[13281] = 8'b10010000;
DRAM[13282] = 8'b10001101;
DRAM[13283] = 8'b10001111;
DRAM[13284] = 8'b10001111;
DRAM[13285] = 8'b10001110;
DRAM[13286] = 8'b10001010;
DRAM[13287] = 8'b10000111;
DRAM[13288] = 8'b10000110;
DRAM[13289] = 8'b10000000;
DRAM[13290] = 8'b01111111;
DRAM[13291] = 8'b01111001;
DRAM[13292] = 8'b01111100;
DRAM[13293] = 8'b10000100;
DRAM[13294] = 8'b01111001;
DRAM[13295] = 8'b10101011;
DRAM[13296] = 8'b11010010;
DRAM[13297] = 8'b11010100;
DRAM[13298] = 8'b11010101;
DRAM[13299] = 8'b11010011;
DRAM[13300] = 8'b11000010;
DRAM[13301] = 8'b10010111;
DRAM[13302] = 8'b01000111;
DRAM[13303] = 8'b01001100;
DRAM[13304] = 8'b01011111;
DRAM[13305] = 8'b01011100;
DRAM[13306] = 8'b01011011;
DRAM[13307] = 8'b01101101;
DRAM[13308] = 8'b01101101;
DRAM[13309] = 8'b01100010;
DRAM[13310] = 8'b01011000;
DRAM[13311] = 8'b01100100;
DRAM[13312] = 8'b01000000;
DRAM[13313] = 8'b01110100;
DRAM[13314] = 8'b10010011;
DRAM[13315] = 8'b10100100;
DRAM[13316] = 8'b10011010;
DRAM[13317] = 8'b01110101;
DRAM[13318] = 8'b00110001;
DRAM[13319] = 8'b01010000;
DRAM[13320] = 8'b10001100;
DRAM[13321] = 8'b10100100;
DRAM[13322] = 8'b10110001;
DRAM[13323] = 8'b10101111;
DRAM[13324] = 8'b10110011;
DRAM[13325] = 8'b10110000;
DRAM[13326] = 8'b10011111;
DRAM[13327] = 8'b10101010;
DRAM[13328] = 8'b01111000;
DRAM[13329] = 8'b01000000;
DRAM[13330] = 8'b00101000;
DRAM[13331] = 8'b00101011;
DRAM[13332] = 8'b00101011;
DRAM[13333] = 8'b00111110;
DRAM[13334] = 8'b00110101;
DRAM[13335] = 8'b00110101;
DRAM[13336] = 8'b00101101;
DRAM[13337] = 8'b00111000;
DRAM[13338] = 8'b01100100;
DRAM[13339] = 8'b01000000;
DRAM[13340] = 8'b00101111;
DRAM[13341] = 8'b01000001;
DRAM[13342] = 8'b01000000;
DRAM[13343] = 8'b00111101;
DRAM[13344] = 8'b01010111;
DRAM[13345] = 8'b01000100;
DRAM[13346] = 8'b01001100;
DRAM[13347] = 8'b01001100;
DRAM[13348] = 8'b01011110;
DRAM[13349] = 8'b01101100;
DRAM[13350] = 8'b01110101;
DRAM[13351] = 8'b10000101;
DRAM[13352] = 8'b10011110;
DRAM[13353] = 8'b01101101;
DRAM[13354] = 8'b01001101;
DRAM[13355] = 8'b01101101;
DRAM[13356] = 8'b10100001;
DRAM[13357] = 8'b00100100;
DRAM[13358] = 8'b00100110;
DRAM[13359] = 8'b01001010;
DRAM[13360] = 8'b00111010;
DRAM[13361] = 8'b00110010;
DRAM[13362] = 8'b00101100;
DRAM[13363] = 8'b00110110;
DRAM[13364] = 8'b00111101;
DRAM[13365] = 8'b00110110;
DRAM[13366] = 8'b00101110;
DRAM[13367] = 8'b01000000;
DRAM[13368] = 8'b01011010;
DRAM[13369] = 8'b01110100;
DRAM[13370] = 8'b01001001;
DRAM[13371] = 8'b00111001;
DRAM[13372] = 8'b01100100;
DRAM[13373] = 8'b01110100;
DRAM[13374] = 8'b10000010;
DRAM[13375] = 8'b10000011;
DRAM[13376] = 8'b10000101;
DRAM[13377] = 8'b10001000;
DRAM[13378] = 8'b10001100;
DRAM[13379] = 8'b10001010;
DRAM[13380] = 8'b10001011;
DRAM[13381] = 8'b10001111;
DRAM[13382] = 8'b10010001;
DRAM[13383] = 8'b10010101;
DRAM[13384] = 8'b10011001;
DRAM[13385] = 8'b10011111;
DRAM[13386] = 8'b10100011;
DRAM[13387] = 8'b10100110;
DRAM[13388] = 8'b10101100;
DRAM[13389] = 8'b10110000;
DRAM[13390] = 8'b10110100;
DRAM[13391] = 8'b10110110;
DRAM[13392] = 8'b10111110;
DRAM[13393] = 8'b11000011;
DRAM[13394] = 8'b11000111;
DRAM[13395] = 8'b11001100;
DRAM[13396] = 8'b11010001;
DRAM[13397] = 8'b11010011;
DRAM[13398] = 8'b11011001;
DRAM[13399] = 8'b11011100;
DRAM[13400] = 8'b01101100;
DRAM[13401] = 8'b00101101;
DRAM[13402] = 8'b00111000;
DRAM[13403] = 8'b00111010;
DRAM[13404] = 8'b00101001;
DRAM[13405] = 8'b10011010;
DRAM[13406] = 8'b10001000;
DRAM[13407] = 8'b10010001;
DRAM[13408] = 8'b10010011;
DRAM[13409] = 8'b10010001;
DRAM[13410] = 8'b10001111;
DRAM[13411] = 8'b10010001;
DRAM[13412] = 8'b10001111;
DRAM[13413] = 8'b10001111;
DRAM[13414] = 8'b10001011;
DRAM[13415] = 8'b10001010;
DRAM[13416] = 8'b10000111;
DRAM[13417] = 8'b10000100;
DRAM[13418] = 8'b10000000;
DRAM[13419] = 8'b01111111;
DRAM[13420] = 8'b10000100;
DRAM[13421] = 8'b10001001;
DRAM[13422] = 8'b10000011;
DRAM[13423] = 8'b11000000;
DRAM[13424] = 8'b11010111;
DRAM[13425] = 8'b11010101;
DRAM[13426] = 8'b11010100;
DRAM[13427] = 8'b11010001;
DRAM[13428] = 8'b10111001;
DRAM[13429] = 8'b01101100;
DRAM[13430] = 8'b01001010;
DRAM[13431] = 8'b01011110;
DRAM[13432] = 8'b01011100;
DRAM[13433] = 8'b01100001;
DRAM[13434] = 8'b01101000;
DRAM[13435] = 8'b01110000;
DRAM[13436] = 8'b01100010;
DRAM[13437] = 8'b01011110;
DRAM[13438] = 8'b01100011;
DRAM[13439] = 8'b01101000;
DRAM[13440] = 8'b00101001;
DRAM[13441] = 8'b01011000;
DRAM[13442] = 8'b10010010;
DRAM[13443] = 8'b10100111;
DRAM[13444] = 8'b10100010;
DRAM[13445] = 8'b10000001;
DRAM[13446] = 8'b00110000;
DRAM[13447] = 8'b01000111;
DRAM[13448] = 8'b10001011;
DRAM[13449] = 8'b10100110;
DRAM[13450] = 8'b10110000;
DRAM[13451] = 8'b10110001;
DRAM[13452] = 8'b10110000;
DRAM[13453] = 8'b10110000;
DRAM[13454] = 8'b10100010;
DRAM[13455] = 8'b10001010;
DRAM[13456] = 8'b10001000;
DRAM[13457] = 8'b01000101;
DRAM[13458] = 8'b00101001;
DRAM[13459] = 8'b00101011;
DRAM[13460] = 8'b00101110;
DRAM[13461] = 8'b01000111;
DRAM[13462] = 8'b00101101;
DRAM[13463] = 8'b00110011;
DRAM[13464] = 8'b00110100;
DRAM[13465] = 8'b01000111;
DRAM[13466] = 8'b01101101;
DRAM[13467] = 8'b00111110;
DRAM[13468] = 8'b00110010;
DRAM[13469] = 8'b00100110;
DRAM[13470] = 8'b01001101;
DRAM[13471] = 8'b00110010;
DRAM[13472] = 8'b01001001;
DRAM[13473] = 8'b01011100;
DRAM[13474] = 8'b01010110;
DRAM[13475] = 8'b01100010;
DRAM[13476] = 8'b01001110;
DRAM[13477] = 8'b01101000;
DRAM[13478] = 8'b01101110;
DRAM[13479] = 8'b01111010;
DRAM[13480] = 8'b10100001;
DRAM[13481] = 8'b01110010;
DRAM[13482] = 8'b00100111;
DRAM[13483] = 8'b01101110;
DRAM[13484] = 8'b11000101;
DRAM[13485] = 8'b00100110;
DRAM[13486] = 8'b00100110;
DRAM[13487] = 8'b01000100;
DRAM[13488] = 8'b01000000;
DRAM[13489] = 8'b00110011;
DRAM[13490] = 8'b00101110;
DRAM[13491] = 8'b00110100;
DRAM[13492] = 8'b01000101;
DRAM[13493] = 8'b00110100;
DRAM[13494] = 8'b00110001;
DRAM[13495] = 8'b00111011;
DRAM[13496] = 8'b01100100;
DRAM[13497] = 8'b01110011;
DRAM[13498] = 8'b01000110;
DRAM[13499] = 8'b00110011;
DRAM[13500] = 8'b01011101;
DRAM[13501] = 8'b01111010;
DRAM[13502] = 8'b10000100;
DRAM[13503] = 8'b10000100;
DRAM[13504] = 8'b10000101;
DRAM[13505] = 8'b10000111;
DRAM[13506] = 8'b10001011;
DRAM[13507] = 8'b10001110;
DRAM[13508] = 8'b10001101;
DRAM[13509] = 8'b10001101;
DRAM[13510] = 8'b10010000;
DRAM[13511] = 8'b10010101;
DRAM[13512] = 8'b10011000;
DRAM[13513] = 8'b10011100;
DRAM[13514] = 8'b10100000;
DRAM[13515] = 8'b10100100;
DRAM[13516] = 8'b10101000;
DRAM[13517] = 8'b10101100;
DRAM[13518] = 8'b10110010;
DRAM[13519] = 8'b10110110;
DRAM[13520] = 8'b10111100;
DRAM[13521] = 8'b11000000;
DRAM[13522] = 8'b11000111;
DRAM[13523] = 8'b11001100;
DRAM[13524] = 8'b11001111;
DRAM[13525] = 8'b11010010;
DRAM[13526] = 8'b11011000;
DRAM[13527] = 8'b11011101;
DRAM[13528] = 8'b11001110;
DRAM[13529] = 8'b00100110;
DRAM[13530] = 8'b00110001;
DRAM[13531] = 8'b00110011;
DRAM[13532] = 8'b00101000;
DRAM[13533] = 8'b10011110;
DRAM[13534] = 8'b10000111;
DRAM[13535] = 8'b10010111;
DRAM[13536] = 8'b10010011;
DRAM[13537] = 8'b10010001;
DRAM[13538] = 8'b10001110;
DRAM[13539] = 8'b10010000;
DRAM[13540] = 8'b10001100;
DRAM[13541] = 8'b10001100;
DRAM[13542] = 8'b10001010;
DRAM[13543] = 8'b10001010;
DRAM[13544] = 8'b10000110;
DRAM[13545] = 8'b10000011;
DRAM[13546] = 8'b10000001;
DRAM[13547] = 8'b01111101;
DRAM[13548] = 8'b10000000;
DRAM[13549] = 8'b10010110;
DRAM[13550] = 8'b10100100;
DRAM[13551] = 8'b11000111;
DRAM[13552] = 8'b11011000;
DRAM[13553] = 8'b11010110;
DRAM[13554] = 8'b11010100;
DRAM[13555] = 8'b11001110;
DRAM[13556] = 8'b10100000;
DRAM[13557] = 8'b01010011;
DRAM[13558] = 8'b01010111;
DRAM[13559] = 8'b01011011;
DRAM[13560] = 8'b01100001;
DRAM[13561] = 8'b01101000;
DRAM[13562] = 8'b01110000;
DRAM[13563] = 8'b01100100;
DRAM[13564] = 8'b01011010;
DRAM[13565] = 8'b01100010;
DRAM[13566] = 8'b01101000;
DRAM[13567] = 8'b01100100;
DRAM[13568] = 8'b00100100;
DRAM[13569] = 8'b01001010;
DRAM[13570] = 8'b10010010;
DRAM[13571] = 8'b10101010;
DRAM[13572] = 8'b10100110;
DRAM[13573] = 8'b10001100;
DRAM[13574] = 8'b00101110;
DRAM[13575] = 8'b01000100;
DRAM[13576] = 8'b10001011;
DRAM[13577] = 8'b10100110;
DRAM[13578] = 8'b10110011;
DRAM[13579] = 8'b10110000;
DRAM[13580] = 8'b10110001;
DRAM[13581] = 8'b10110010;
DRAM[13582] = 8'b10100100;
DRAM[13583] = 8'b10001010;
DRAM[13584] = 8'b01101011;
DRAM[13585] = 8'b01010011;
DRAM[13586] = 8'b00110000;
DRAM[13587] = 8'b00101011;
DRAM[13588] = 8'b00111000;
DRAM[13589] = 8'b00110001;
DRAM[13590] = 8'b00101100;
DRAM[13591] = 8'b00110001;
DRAM[13592] = 8'b00101010;
DRAM[13593] = 8'b01001000;
DRAM[13594] = 8'b01011110;
DRAM[13595] = 8'b00110100;
DRAM[13596] = 8'b00111100;
DRAM[13597] = 8'b00101011;
DRAM[13598] = 8'b00110001;
DRAM[13599] = 8'b01001111;
DRAM[13600] = 8'b01010011;
DRAM[13601] = 8'b00111100;
DRAM[13602] = 8'b01010101;
DRAM[13603] = 8'b01101110;
DRAM[13604] = 8'b01011101;
DRAM[13605] = 8'b01010100;
DRAM[13606] = 8'b01100111;
DRAM[13607] = 8'b10010110;
DRAM[13608] = 8'b10001100;
DRAM[13609] = 8'b01010110;
DRAM[13610] = 8'b00111001;
DRAM[13611] = 8'b10000001;
DRAM[13612] = 8'b10111000;
DRAM[13613] = 8'b00101000;
DRAM[13614] = 8'b00100100;
DRAM[13615] = 8'b01000000;
DRAM[13616] = 8'b01010001;
DRAM[13617] = 8'b00110010;
DRAM[13618] = 8'b00101111;
DRAM[13619] = 8'b00110101;
DRAM[13620] = 8'b00111111;
DRAM[13621] = 8'b00110000;
DRAM[13622] = 8'b00110001;
DRAM[13623] = 8'b00111111;
DRAM[13624] = 8'b01101010;
DRAM[13625] = 8'b01101011;
DRAM[13626] = 8'b01010010;
DRAM[13627] = 8'b00110001;
DRAM[13628] = 8'b01101000;
DRAM[13629] = 8'b01111001;
DRAM[13630] = 8'b10000010;
DRAM[13631] = 8'b10000000;
DRAM[13632] = 8'b10000111;
DRAM[13633] = 8'b10000110;
DRAM[13634] = 8'b10001001;
DRAM[13635] = 8'b10001010;
DRAM[13636] = 8'b10001100;
DRAM[13637] = 8'b10001101;
DRAM[13638] = 8'b10010100;
DRAM[13639] = 8'b10010101;
DRAM[13640] = 8'b10010110;
DRAM[13641] = 8'b10011010;
DRAM[13642] = 8'b10011101;
DRAM[13643] = 8'b10100011;
DRAM[13644] = 8'b10100111;
DRAM[13645] = 8'b10101101;
DRAM[13646] = 8'b10110001;
DRAM[13647] = 8'b10110110;
DRAM[13648] = 8'b10111001;
DRAM[13649] = 8'b10111110;
DRAM[13650] = 8'b11000110;
DRAM[13651] = 8'b11001011;
DRAM[13652] = 8'b11010000;
DRAM[13653] = 8'b11010010;
DRAM[13654] = 8'b11010111;
DRAM[13655] = 8'b11011010;
DRAM[13656] = 8'b11011101;
DRAM[13657] = 8'b01110011;
DRAM[13658] = 8'b00101010;
DRAM[13659] = 8'b00101000;
DRAM[13660] = 8'b00111000;
DRAM[13661] = 8'b10011010;
DRAM[13662] = 8'b10001011;
DRAM[13663] = 8'b10010101;
DRAM[13664] = 8'b10010101;
DRAM[13665] = 8'b10010010;
DRAM[13666] = 8'b10010000;
DRAM[13667] = 8'b10001110;
DRAM[13668] = 8'b10001110;
DRAM[13669] = 8'b10001001;
DRAM[13670] = 8'b10001000;
DRAM[13671] = 8'b10000110;
DRAM[13672] = 8'b10000101;
DRAM[13673] = 8'b10000001;
DRAM[13674] = 8'b01111100;
DRAM[13675] = 8'b01111001;
DRAM[13676] = 8'b10011001;
DRAM[13677] = 8'b10111000;
DRAM[13678] = 8'b11000011;
DRAM[13679] = 8'b11010001;
DRAM[13680] = 8'b11010111;
DRAM[13681] = 8'b11010110;
DRAM[13682] = 8'b11010011;
DRAM[13683] = 8'b11000100;
DRAM[13684] = 8'b01111100;
DRAM[13685] = 8'b01010111;
DRAM[13686] = 8'b01011101;
DRAM[13687] = 8'b01011111;
DRAM[13688] = 8'b01100110;
DRAM[13689] = 8'b01101111;
DRAM[13690] = 8'b01101001;
DRAM[13691] = 8'b01011010;
DRAM[13692] = 8'b01011010;
DRAM[13693] = 8'b01100100;
DRAM[13694] = 8'b01100011;
DRAM[13695] = 8'b01100110;
DRAM[13696] = 8'b00100110;
DRAM[13697] = 8'b00111001;
DRAM[13698] = 8'b10000110;
DRAM[13699] = 8'b10101001;
DRAM[13700] = 8'b10100111;
DRAM[13701] = 8'b10000011;
DRAM[13702] = 8'b00101100;
DRAM[13703] = 8'b01000010;
DRAM[13704] = 8'b10000111;
DRAM[13705] = 8'b10100110;
DRAM[13706] = 8'b10110011;
DRAM[13707] = 8'b10110000;
DRAM[13708] = 8'b10110011;
DRAM[13709] = 8'b10110100;
DRAM[13710] = 8'b10100100;
DRAM[13711] = 8'b10001100;
DRAM[13712] = 8'b10010110;
DRAM[13713] = 8'b00101101;
DRAM[13714] = 8'b00110001;
DRAM[13715] = 8'b00110100;
DRAM[13716] = 8'b00110100;
DRAM[13717] = 8'b00110001;
DRAM[13718] = 8'b00101011;
DRAM[13719] = 8'b00110011;
DRAM[13720] = 8'b00101100;
DRAM[13721] = 8'b01101001;
DRAM[13722] = 8'b01011001;
DRAM[13723] = 8'b00101000;
DRAM[13724] = 8'b01000100;
DRAM[13725] = 8'b00110111;
DRAM[13726] = 8'b00110000;
DRAM[13727] = 8'b00111000;
DRAM[13728] = 8'b00110010;
DRAM[13729] = 8'b01000101;
DRAM[13730] = 8'b01001001;
DRAM[13731] = 8'b01100011;
DRAM[13732] = 8'b01100010;
DRAM[13733] = 8'b01001111;
DRAM[13734] = 8'b01100110;
DRAM[13735] = 8'b10001100;
DRAM[13736] = 8'b10010011;
DRAM[13737] = 8'b01101101;
DRAM[13738] = 8'b00101010;
DRAM[13739] = 8'b10000000;
DRAM[13740] = 8'b10000101;
DRAM[13741] = 8'b00101010;
DRAM[13742] = 8'b00101100;
DRAM[13743] = 8'b01000000;
DRAM[13744] = 8'b01001011;
DRAM[13745] = 8'b00111000;
DRAM[13746] = 8'b00110010;
DRAM[13747] = 8'b00110110;
DRAM[13748] = 8'b00111110;
DRAM[13749] = 8'b00101100;
DRAM[13750] = 8'b00110100;
DRAM[13751] = 8'b01001000;
DRAM[13752] = 8'b01100110;
DRAM[13753] = 8'b01101111;
DRAM[13754] = 8'b01011100;
DRAM[13755] = 8'b00110100;
DRAM[13756] = 8'b01100011;
DRAM[13757] = 8'b01111101;
DRAM[13758] = 8'b10000001;
DRAM[13759] = 8'b10000011;
DRAM[13760] = 8'b10001001;
DRAM[13761] = 8'b10001001;
DRAM[13762] = 8'b10001001;
DRAM[13763] = 8'b10001000;
DRAM[13764] = 8'b10001011;
DRAM[13765] = 8'b10001101;
DRAM[13766] = 8'b10001111;
DRAM[13767] = 8'b10010001;
DRAM[13768] = 8'b10010101;
DRAM[13769] = 8'b10011011;
DRAM[13770] = 8'b10011100;
DRAM[13771] = 8'b10100000;
DRAM[13772] = 8'b10100111;
DRAM[13773] = 8'b10101001;
DRAM[13774] = 8'b10101111;
DRAM[13775] = 8'b10110100;
DRAM[13776] = 8'b10111011;
DRAM[13777] = 8'b10111101;
DRAM[13778] = 8'b11000101;
DRAM[13779] = 8'b11001011;
DRAM[13780] = 8'b11010000;
DRAM[13781] = 8'b11010011;
DRAM[13782] = 8'b11010101;
DRAM[13783] = 8'b11011000;
DRAM[13784] = 8'b11011100;
DRAM[13785] = 8'b11001001;
DRAM[13786] = 8'b00100000;
DRAM[13787] = 8'b00100101;
DRAM[13788] = 8'b01010010;
DRAM[13789] = 8'b10010001;
DRAM[13790] = 8'b10010001;
DRAM[13791] = 8'b10010101;
DRAM[13792] = 8'b10010010;
DRAM[13793] = 8'b10010000;
DRAM[13794] = 8'b10010011;
DRAM[13795] = 8'b10001101;
DRAM[13796] = 8'b10001101;
DRAM[13797] = 8'b10001010;
DRAM[13798] = 8'b10000111;
DRAM[13799] = 8'b10000101;
DRAM[13800] = 8'b10000100;
DRAM[13801] = 8'b01111111;
DRAM[13802] = 8'b01111001;
DRAM[13803] = 8'b10001110;
DRAM[13804] = 8'b10111111;
DRAM[13805] = 8'b11001011;
DRAM[13806] = 8'b11001010;
DRAM[13807] = 8'b11010101;
DRAM[13808] = 8'b11011001;
DRAM[13809] = 8'b11010111;
DRAM[13810] = 8'b11001110;
DRAM[13811] = 8'b10101000;
DRAM[13812] = 8'b01100010;
DRAM[13813] = 8'b01011010;
DRAM[13814] = 8'b01011100;
DRAM[13815] = 8'b01100111;
DRAM[13816] = 8'b01101111;
DRAM[13817] = 8'b01110010;
DRAM[13818] = 8'b01011110;
DRAM[13819] = 8'b01011011;
DRAM[13820] = 8'b01100100;
DRAM[13821] = 8'b01100110;
DRAM[13822] = 8'b01100000;
DRAM[13823] = 8'b01101000;
DRAM[13824] = 8'b00011110;
DRAM[13825] = 8'b00101111;
DRAM[13826] = 8'b10000100;
DRAM[13827] = 8'b10100100;
DRAM[13828] = 8'b10101000;
DRAM[13829] = 8'b10000101;
DRAM[13830] = 8'b00101011;
DRAM[13831] = 8'b00111111;
DRAM[13832] = 8'b10001010;
DRAM[13833] = 8'b10100110;
DRAM[13834] = 8'b10110010;
DRAM[13835] = 8'b10110010;
DRAM[13836] = 8'b10110010;
DRAM[13837] = 8'b10110011;
DRAM[13838] = 8'b10100100;
DRAM[13839] = 8'b10001100;
DRAM[13840] = 8'b01111101;
DRAM[13841] = 8'b00110101;
DRAM[13842] = 8'b00110100;
DRAM[13843] = 8'b00110111;
DRAM[13844] = 8'b00101101;
DRAM[13845] = 8'b00101101;
DRAM[13846] = 8'b00101110;
DRAM[13847] = 8'b00101000;
DRAM[13848] = 8'b00110101;
DRAM[13849] = 8'b10001100;
DRAM[13850] = 8'b01001110;
DRAM[13851] = 8'b00101110;
DRAM[13852] = 8'b00110100;
DRAM[13853] = 8'b00111011;
DRAM[13854] = 8'b00110100;
DRAM[13855] = 8'b00110011;
DRAM[13856] = 8'b00110010;
DRAM[13857] = 8'b00110000;
DRAM[13858] = 8'b01001001;
DRAM[13859] = 8'b01011010;
DRAM[13860] = 8'b01101010;
DRAM[13861] = 8'b01000000;
DRAM[13862] = 8'b01100010;
DRAM[13863] = 8'b10001101;
DRAM[13864] = 8'b10011001;
DRAM[13865] = 8'b01110100;
DRAM[13866] = 8'b01101100;
DRAM[13867] = 8'b10001110;
DRAM[13868] = 8'b10001111;
DRAM[13869] = 8'b01101001;
DRAM[13870] = 8'b00110111;
DRAM[13871] = 8'b00111011;
DRAM[13872] = 8'b01000101;
DRAM[13873] = 8'b00110101;
DRAM[13874] = 8'b00111001;
DRAM[13875] = 8'b00110011;
DRAM[13876] = 8'b00110010;
DRAM[13877] = 8'b00111000;
DRAM[13878] = 8'b00111010;
DRAM[13879] = 8'b01011011;
DRAM[13880] = 8'b01111000;
DRAM[13881] = 8'b01111010;
DRAM[13882] = 8'b01100100;
DRAM[13883] = 8'b00111111;
DRAM[13884] = 8'b01101000;
DRAM[13885] = 8'b01111111;
DRAM[13886] = 8'b10000100;
DRAM[13887] = 8'b10000110;
DRAM[13888] = 8'b10001100;
DRAM[13889] = 8'b10001000;
DRAM[13890] = 8'b10001001;
DRAM[13891] = 8'b10001010;
DRAM[13892] = 8'b10001010;
DRAM[13893] = 8'b10001011;
DRAM[13894] = 8'b10010010;
DRAM[13895] = 8'b10010001;
DRAM[13896] = 8'b10010011;
DRAM[13897] = 8'b10011000;
DRAM[13898] = 8'b10011011;
DRAM[13899] = 8'b10011111;
DRAM[13900] = 8'b10100011;
DRAM[13901] = 8'b10100111;
DRAM[13902] = 8'b10101111;
DRAM[13903] = 8'b10110010;
DRAM[13904] = 8'b10111001;
DRAM[13905] = 8'b10111101;
DRAM[13906] = 8'b11000100;
DRAM[13907] = 8'b11001011;
DRAM[13908] = 8'b11010000;
DRAM[13909] = 8'b11010011;
DRAM[13910] = 8'b11010101;
DRAM[13911] = 8'b11010111;
DRAM[13912] = 8'b11011011;
DRAM[13913] = 8'b11011101;
DRAM[13914] = 8'b01001000;
DRAM[13915] = 8'b00011111;
DRAM[13916] = 8'b01100000;
DRAM[13917] = 8'b10010001;
DRAM[13918] = 8'b10010101;
DRAM[13919] = 8'b10010100;
DRAM[13920] = 8'b10010010;
DRAM[13921] = 8'b10010010;
DRAM[13922] = 8'b10010000;
DRAM[13923] = 8'b10001111;
DRAM[13924] = 8'b10001011;
DRAM[13925] = 8'b10001010;
DRAM[13926] = 8'b10000101;
DRAM[13927] = 8'b10000010;
DRAM[13928] = 8'b10000000;
DRAM[13929] = 8'b01111110;
DRAM[13930] = 8'b01111001;
DRAM[13931] = 8'b10101010;
DRAM[13932] = 8'b11010100;
DRAM[13933] = 8'b11010110;
DRAM[13934] = 8'b11001101;
DRAM[13935] = 8'b11010110;
DRAM[13936] = 8'b11011001;
DRAM[13937] = 8'b11010100;
DRAM[13938] = 8'b11000011;
DRAM[13939] = 8'b10000110;
DRAM[13940] = 8'b01100000;
DRAM[13941] = 8'b01011100;
DRAM[13942] = 8'b01011100;
DRAM[13943] = 8'b01101011;
DRAM[13944] = 8'b01110010;
DRAM[13945] = 8'b01101101;
DRAM[13946] = 8'b01011100;
DRAM[13947] = 8'b01011011;
DRAM[13948] = 8'b01100111;
DRAM[13949] = 8'b01100111;
DRAM[13950] = 8'b01100101;
DRAM[13951] = 8'b01100001;
DRAM[13952] = 8'b00011111;
DRAM[13953] = 8'b00101011;
DRAM[13954] = 8'b01111100;
DRAM[13955] = 8'b10100111;
DRAM[13956] = 8'b10101011;
DRAM[13957] = 8'b10001010;
DRAM[13958] = 8'b00110100;
DRAM[13959] = 8'b00111101;
DRAM[13960] = 8'b10001000;
DRAM[13961] = 8'b10100110;
DRAM[13962] = 8'b10110010;
DRAM[13963] = 8'b10110000;
DRAM[13964] = 8'b10110100;
DRAM[13965] = 8'b10110011;
DRAM[13966] = 8'b10100101;
DRAM[13967] = 8'b10001111;
DRAM[13968] = 8'b01100000;
DRAM[13969] = 8'b00111010;
DRAM[13970] = 8'b00110101;
DRAM[13971] = 8'b00101001;
DRAM[13972] = 8'b00101011;
DRAM[13973] = 8'b00101110;
DRAM[13974] = 8'b00101110;
DRAM[13975] = 8'b00101110;
DRAM[13976] = 8'b01100101;
DRAM[13977] = 8'b01011000;
DRAM[13978] = 8'b00111110;
DRAM[13979] = 8'b00101101;
DRAM[13980] = 8'b00110101;
DRAM[13981] = 8'b01000100;
DRAM[13982] = 8'b00110001;
DRAM[13983] = 8'b00100101;
DRAM[13984] = 8'b00111101;
DRAM[13985] = 8'b00101011;
DRAM[13986] = 8'b01000101;
DRAM[13987] = 8'b01000101;
DRAM[13988] = 8'b01110011;
DRAM[13989] = 8'b01011001;
DRAM[13990] = 8'b01110111;
DRAM[13991] = 8'b10001010;
DRAM[13992] = 8'b01110011;
DRAM[13993] = 8'b10000001;
DRAM[13994] = 8'b10001111;
DRAM[13995] = 8'b10010101;
DRAM[13996] = 8'b00111001;
DRAM[13997] = 8'b00111000;
DRAM[13998] = 8'b00111010;
DRAM[13999] = 8'b00110100;
DRAM[14000] = 8'b01000001;
DRAM[14001] = 8'b00111000;
DRAM[14002] = 8'b00110111;
DRAM[14003] = 8'b00110111;
DRAM[14004] = 8'b00110010;
DRAM[14005] = 8'b00110111;
DRAM[14006] = 8'b01001000;
DRAM[14007] = 8'b01110011;
DRAM[14008] = 8'b01111100;
DRAM[14009] = 8'b01111010;
DRAM[14010] = 8'b01010110;
DRAM[14011] = 8'b01000010;
DRAM[14012] = 8'b01100110;
DRAM[14013] = 8'b01111100;
DRAM[14014] = 8'b10000010;
DRAM[14015] = 8'b10000101;
DRAM[14016] = 8'b10001011;
DRAM[14017] = 8'b10001010;
DRAM[14018] = 8'b10001000;
DRAM[14019] = 8'b10001000;
DRAM[14020] = 8'b10001011;
DRAM[14021] = 8'b10001100;
DRAM[14022] = 8'b10001110;
DRAM[14023] = 8'b10010000;
DRAM[14024] = 8'b10010010;
DRAM[14025] = 8'b10010101;
DRAM[14026] = 8'b10011011;
DRAM[14027] = 8'b10011110;
DRAM[14028] = 8'b10100000;
DRAM[14029] = 8'b10100101;
DRAM[14030] = 8'b10101110;
DRAM[14031] = 8'b10110001;
DRAM[14032] = 8'b10110101;
DRAM[14033] = 8'b10111101;
DRAM[14034] = 8'b11000010;
DRAM[14035] = 8'b11001001;
DRAM[14036] = 8'b11001101;
DRAM[14037] = 8'b11001111;
DRAM[14038] = 8'b11010011;
DRAM[14039] = 8'b11010101;
DRAM[14040] = 8'b11011000;
DRAM[14041] = 8'b11011101;
DRAM[14042] = 8'b01111010;
DRAM[14043] = 8'b00011111;
DRAM[14044] = 8'b01011111;
DRAM[14045] = 8'b10001111;
DRAM[14046] = 8'b10010101;
DRAM[14047] = 8'b10010000;
DRAM[14048] = 8'b10010010;
DRAM[14049] = 8'b10010000;
DRAM[14050] = 8'b10001101;
DRAM[14051] = 8'b10001101;
DRAM[14052] = 8'b10001101;
DRAM[14053] = 8'b10001010;
DRAM[14054] = 8'b10000101;
DRAM[14055] = 8'b10000100;
DRAM[14056] = 8'b01111111;
DRAM[14057] = 8'b01111010;
DRAM[14058] = 8'b01111011;
DRAM[14059] = 8'b10111101;
DRAM[14060] = 8'b11011000;
DRAM[14061] = 8'b11010100;
DRAM[14062] = 8'b11010001;
DRAM[14063] = 8'b11010111;
DRAM[14064] = 8'b11011000;
DRAM[14065] = 8'b11010001;
DRAM[14066] = 8'b10101011;
DRAM[14067] = 8'b01110101;
DRAM[14068] = 8'b01100110;
DRAM[14069] = 8'b01011111;
DRAM[14070] = 8'b01011110;
DRAM[14071] = 8'b01110000;
DRAM[14072] = 8'b01110000;
DRAM[14073] = 8'b01100011;
DRAM[14074] = 8'b01011010;
DRAM[14075] = 8'b01100011;
DRAM[14076] = 8'b01101001;
DRAM[14077] = 8'b01100010;
DRAM[14078] = 8'b01100000;
DRAM[14079] = 8'b01010011;
DRAM[14080] = 8'b00011111;
DRAM[14081] = 8'b00101000;
DRAM[14082] = 8'b01111111;
DRAM[14083] = 8'b10100011;
DRAM[14084] = 8'b10101001;
DRAM[14085] = 8'b10001100;
DRAM[14086] = 8'b01000010;
DRAM[14087] = 8'b00111000;
DRAM[14088] = 8'b10001000;
DRAM[14089] = 8'b10100111;
DRAM[14090] = 8'b10110001;
DRAM[14091] = 8'b10101110;
DRAM[14092] = 8'b10101011;
DRAM[14093] = 8'b10101110;
DRAM[14094] = 8'b10100010;
DRAM[14095] = 8'b10010000;
DRAM[14096] = 8'b01111000;
DRAM[14097] = 8'b00111000;
DRAM[14098] = 8'b00101111;
DRAM[14099] = 8'b00110000;
DRAM[14100] = 8'b00101110;
DRAM[14101] = 8'b00110010;
DRAM[14102] = 8'b00111111;
DRAM[14103] = 8'b01000010;
DRAM[14104] = 8'b00101110;
DRAM[14105] = 8'b01001111;
DRAM[14106] = 8'b01001110;
DRAM[14107] = 8'b00101100;
DRAM[14108] = 8'b00110110;
DRAM[14109] = 8'b00111010;
DRAM[14110] = 8'b00101010;
DRAM[14111] = 8'b00101110;
DRAM[14112] = 8'b01000000;
DRAM[14113] = 8'b00101111;
DRAM[14114] = 8'b01010100;
DRAM[14115] = 8'b00110011;
DRAM[14116] = 8'b00110101;
DRAM[14117] = 8'b01110001;
DRAM[14118] = 8'b10000100;
DRAM[14119] = 8'b10000110;
DRAM[14120] = 8'b01101111;
DRAM[14121] = 8'b01010001;
DRAM[14122] = 8'b01111000;
DRAM[14123] = 8'b10010010;
DRAM[14124] = 8'b10000011;
DRAM[14125] = 8'b01100100;
DRAM[14126] = 8'b01011010;
DRAM[14127] = 8'b00111010;
DRAM[14128] = 8'b00110111;
DRAM[14129] = 8'b01001000;
DRAM[14130] = 8'b00111010;
DRAM[14131] = 8'b00111010;
DRAM[14132] = 8'b00110000;
DRAM[14133] = 8'b00111101;
DRAM[14134] = 8'b01010010;
DRAM[14135] = 8'b01110111;
DRAM[14136] = 8'b01111110;
DRAM[14137] = 8'b01111100;
DRAM[14138] = 8'b01001110;
DRAM[14139] = 8'b01000111;
DRAM[14140] = 8'b01101110;
DRAM[14141] = 8'b01111110;
DRAM[14142] = 8'b10000101;
DRAM[14143] = 8'b10000111;
DRAM[14144] = 8'b10001011;
DRAM[14145] = 8'b10001110;
DRAM[14146] = 8'b10000111;
DRAM[14147] = 8'b10001001;
DRAM[14148] = 8'b10000111;
DRAM[14149] = 8'b10001010;
DRAM[14150] = 8'b10001100;
DRAM[14151] = 8'b10001110;
DRAM[14152] = 8'b10010001;
DRAM[14153] = 8'b10010100;
DRAM[14154] = 8'b10011000;
DRAM[14155] = 8'b10011101;
DRAM[14156] = 8'b10100001;
DRAM[14157] = 8'b10100101;
DRAM[14158] = 8'b10101001;
DRAM[14159] = 8'b10101110;
DRAM[14160] = 8'b10110110;
DRAM[14161] = 8'b10111100;
DRAM[14162] = 8'b11000000;
DRAM[14163] = 8'b11000111;
DRAM[14164] = 8'b11001100;
DRAM[14165] = 8'b11001110;
DRAM[14166] = 8'b11010010;
DRAM[14167] = 8'b11010100;
DRAM[14168] = 8'b11011000;
DRAM[14169] = 8'b11011011;
DRAM[14170] = 8'b11000001;
DRAM[14171] = 8'b00011001;
DRAM[14172] = 8'b01101100;
DRAM[14173] = 8'b10010000;
DRAM[14174] = 8'b10010011;
DRAM[14175] = 8'b10010001;
DRAM[14176] = 8'b10001101;
DRAM[14177] = 8'b10001101;
DRAM[14178] = 8'b10001010;
DRAM[14179] = 8'b10001011;
DRAM[14180] = 8'b10001011;
DRAM[14181] = 8'b10001001;
DRAM[14182] = 8'b10001000;
DRAM[14183] = 8'b10000110;
DRAM[14184] = 8'b10000000;
DRAM[14185] = 8'b01111100;
DRAM[14186] = 8'b10000011;
DRAM[14187] = 8'b11000100;
DRAM[14188] = 8'b11010110;
DRAM[14189] = 8'b11001111;
DRAM[14190] = 8'b11010001;
DRAM[14191] = 8'b11011001;
DRAM[14192] = 8'b11010110;
DRAM[14193] = 8'b11000101;
DRAM[14194] = 8'b10001110;
DRAM[14195] = 8'b01110111;
DRAM[14196] = 8'b01101001;
DRAM[14197] = 8'b01100010;
DRAM[14198] = 8'b01100101;
DRAM[14199] = 8'b01101100;
DRAM[14200] = 8'b01101100;
DRAM[14201] = 8'b01100001;
DRAM[14202] = 8'b01011011;
DRAM[14203] = 8'b01100110;
DRAM[14204] = 8'b01100111;
DRAM[14205] = 8'b01100010;
DRAM[14206] = 8'b01011000;
DRAM[14207] = 8'b01010010;
DRAM[14208] = 8'b00100000;
DRAM[14209] = 8'b00100111;
DRAM[14210] = 8'b01101000;
DRAM[14211] = 8'b10100011;
DRAM[14212] = 8'b10101100;
DRAM[14213] = 8'b10010100;
DRAM[14214] = 8'b00111110;
DRAM[14215] = 8'b00111001;
DRAM[14216] = 8'b10000110;
DRAM[14217] = 8'b10100110;
DRAM[14218] = 8'b10110001;
DRAM[14219] = 8'b10110001;
DRAM[14220] = 8'b10110000;
DRAM[14221] = 8'b10110001;
DRAM[14222] = 8'b10100100;
DRAM[14223] = 8'b10010100;
DRAM[14224] = 8'b01110011;
DRAM[14225] = 8'b00110100;
DRAM[14226] = 8'b00110000;
DRAM[14227] = 8'b00101110;
DRAM[14228] = 8'b00101111;
DRAM[14229] = 8'b00110000;
DRAM[14230] = 8'b00111000;
DRAM[14231] = 8'b00110101;
DRAM[14232] = 8'b00110100;
DRAM[14233] = 8'b01000001;
DRAM[14234] = 8'b01000100;
DRAM[14235] = 8'b00110011;
DRAM[14236] = 8'b00111100;
DRAM[14237] = 8'b00111000;
DRAM[14238] = 8'b00110000;
DRAM[14239] = 8'b00101110;
DRAM[14240] = 8'b00111101;
DRAM[14241] = 8'b00101111;
DRAM[14242] = 8'b01001111;
DRAM[14243] = 8'b00110101;
DRAM[14244] = 8'b00101111;
DRAM[14245] = 8'b01101100;
DRAM[14246] = 8'b01110100;
DRAM[14247] = 8'b01110110;
DRAM[14248] = 8'b01111000;
DRAM[14249] = 8'b01001011;
DRAM[14250] = 8'b00110100;
DRAM[14251] = 8'b00101010;
DRAM[14252] = 8'b00111011;
DRAM[14253] = 8'b00101010;
DRAM[14254] = 8'b01100100;
DRAM[14255] = 8'b01110100;
DRAM[14256] = 8'b01100100;
DRAM[14257] = 8'b01001100;
DRAM[14258] = 8'b00110101;
DRAM[14259] = 8'b00110100;
DRAM[14260] = 8'b00110010;
DRAM[14261] = 8'b01000111;
DRAM[14262] = 8'b01100010;
DRAM[14263] = 8'b01111100;
DRAM[14264] = 8'b01111111;
DRAM[14265] = 8'b01111111;
DRAM[14266] = 8'b01000001;
DRAM[14267] = 8'b01010111;
DRAM[14268] = 8'b01110101;
DRAM[14269] = 8'b10000100;
DRAM[14270] = 8'b10000110;
DRAM[14271] = 8'b10000111;
DRAM[14272] = 8'b10001010;
DRAM[14273] = 8'b10001100;
DRAM[14274] = 8'b10001010;
DRAM[14275] = 8'b10001010;
DRAM[14276] = 8'b10000111;
DRAM[14277] = 8'b10000111;
DRAM[14278] = 8'b10001011;
DRAM[14279] = 8'b10001101;
DRAM[14280] = 8'b10001110;
DRAM[14281] = 8'b10010101;
DRAM[14282] = 8'b10010111;
DRAM[14283] = 8'b10011010;
DRAM[14284] = 8'b10011110;
DRAM[14285] = 8'b10100001;
DRAM[14286] = 8'b10100111;
DRAM[14287] = 8'b10101000;
DRAM[14288] = 8'b10110001;
DRAM[14289] = 8'b10110111;
DRAM[14290] = 8'b11000010;
DRAM[14291] = 8'b11000100;
DRAM[14292] = 8'b11001000;
DRAM[14293] = 8'b11001101;
DRAM[14294] = 8'b11010000;
DRAM[14295] = 8'b11010100;
DRAM[14296] = 8'b11010101;
DRAM[14297] = 8'b11011000;
DRAM[14298] = 8'b11011001;
DRAM[14299] = 8'b00100110;
DRAM[14300] = 8'b10000001;
DRAM[14301] = 8'b10010000;
DRAM[14302] = 8'b10010001;
DRAM[14303] = 8'b10010100;
DRAM[14304] = 8'b10001111;
DRAM[14305] = 8'b10001110;
DRAM[14306] = 8'b10001011;
DRAM[14307] = 8'b10001010;
DRAM[14308] = 8'b10001010;
DRAM[14309] = 8'b10001010;
DRAM[14310] = 8'b10000110;
DRAM[14311] = 8'b10000100;
DRAM[14312] = 8'b01111110;
DRAM[14313] = 8'b01111100;
DRAM[14314] = 8'b10000111;
DRAM[14315] = 8'b11000111;
DRAM[14316] = 8'b11010111;
DRAM[14317] = 8'b11001011;
DRAM[14318] = 8'b11010000;
DRAM[14319] = 8'b11011010;
DRAM[14320] = 8'b11010010;
DRAM[14321] = 8'b10110001;
DRAM[14322] = 8'b01111110;
DRAM[14323] = 8'b01110100;
DRAM[14324] = 8'b01100111;
DRAM[14325] = 8'b01100001;
DRAM[14326] = 8'b01100110;
DRAM[14327] = 8'b01101001;
DRAM[14328] = 8'b01100011;
DRAM[14329] = 8'b01011000;
DRAM[14330] = 8'b01011110;
DRAM[14331] = 8'b01101000;
DRAM[14332] = 8'b01100010;
DRAM[14333] = 8'b01011100;
DRAM[14334] = 8'b01011011;
DRAM[14335] = 8'b01011001;
DRAM[14336] = 8'b00100011;
DRAM[14337] = 8'b00100100;
DRAM[14338] = 8'b01011101;
DRAM[14339] = 8'b10011110;
DRAM[14340] = 8'b10101011;
DRAM[14341] = 8'b10010011;
DRAM[14342] = 8'b01000010;
DRAM[14343] = 8'b00111110;
DRAM[14344] = 8'b10000101;
DRAM[14345] = 8'b10100100;
DRAM[14346] = 8'b10110000;
DRAM[14347] = 8'b10110001;
DRAM[14348] = 8'b10110010;
DRAM[14349] = 8'b10110011;
DRAM[14350] = 8'b10100100;
DRAM[14351] = 8'b10010011;
DRAM[14352] = 8'b01110001;
DRAM[14353] = 8'b00110101;
DRAM[14354] = 8'b00110100;
DRAM[14355] = 8'b00101010;
DRAM[14356] = 8'b00101011;
DRAM[14357] = 8'b00110000;
DRAM[14358] = 8'b00110101;
DRAM[14359] = 8'b01000000;
DRAM[14360] = 8'b00110000;
DRAM[14361] = 8'b01000001;
DRAM[14362] = 8'b00111111;
DRAM[14363] = 8'b00110111;
DRAM[14364] = 8'b00110000;
DRAM[14365] = 8'b00110110;
DRAM[14366] = 8'b00111110;
DRAM[14367] = 8'b00101000;
DRAM[14368] = 8'b00110101;
DRAM[14369] = 8'b00111011;
DRAM[14370] = 8'b01010101;
DRAM[14371] = 8'b00111011;
DRAM[14372] = 8'b01011010;
DRAM[14373] = 8'b01010110;
DRAM[14374] = 8'b01110101;
DRAM[14375] = 8'b01101011;
DRAM[14376] = 8'b01101011;
DRAM[14377] = 8'b10001011;
DRAM[14378] = 8'b00111001;
DRAM[14379] = 8'b01010000;
DRAM[14380] = 8'b00110000;
DRAM[14381] = 8'b00110111;
DRAM[14382] = 8'b00111011;
DRAM[14383] = 8'b00111001;
DRAM[14384] = 8'b00111001;
DRAM[14385] = 8'b01000110;
DRAM[14386] = 8'b00111001;
DRAM[14387] = 8'b00101100;
DRAM[14388] = 8'b00111101;
DRAM[14389] = 8'b01010010;
DRAM[14390] = 8'b01101001;
DRAM[14391] = 8'b01111100;
DRAM[14392] = 8'b10000010;
DRAM[14393] = 8'b01111001;
DRAM[14394] = 8'b01000001;
DRAM[14395] = 8'b01100001;
DRAM[14396] = 8'b01111111;
DRAM[14397] = 8'b10000101;
DRAM[14398] = 8'b10001001;
DRAM[14399] = 8'b10001011;
DRAM[14400] = 8'b10001101;
DRAM[14401] = 8'b10001101;
DRAM[14402] = 8'b10001101;
DRAM[14403] = 8'b10001000;
DRAM[14404] = 8'b10001000;
DRAM[14405] = 8'b10001000;
DRAM[14406] = 8'b10001011;
DRAM[14407] = 8'b10001011;
DRAM[14408] = 8'b10001101;
DRAM[14409] = 8'b10010011;
DRAM[14410] = 8'b10010100;
DRAM[14411] = 8'b10011100;
DRAM[14412] = 8'b10011110;
DRAM[14413] = 8'b10100010;
DRAM[14414] = 8'b10100110;
DRAM[14415] = 8'b10101000;
DRAM[14416] = 8'b10101110;
DRAM[14417] = 8'b10111000;
DRAM[14418] = 8'b10111111;
DRAM[14419] = 8'b11000110;
DRAM[14420] = 8'b11000111;
DRAM[14421] = 8'b11001101;
DRAM[14422] = 8'b11001111;
DRAM[14423] = 8'b11010010;
DRAM[14424] = 8'b11010101;
DRAM[14425] = 8'b11010101;
DRAM[14426] = 8'b11011000;
DRAM[14427] = 8'b01101100;
DRAM[14428] = 8'b10001010;
DRAM[14429] = 8'b10010001;
DRAM[14430] = 8'b10010111;
DRAM[14431] = 8'b10010010;
DRAM[14432] = 8'b10001101;
DRAM[14433] = 8'b10001110;
DRAM[14434] = 8'b10001101;
DRAM[14435] = 8'b10001101;
DRAM[14436] = 8'b10001101;
DRAM[14437] = 8'b10001011;
DRAM[14438] = 8'b10001000;
DRAM[14439] = 8'b10000011;
DRAM[14440] = 8'b10000000;
DRAM[14441] = 8'b10000011;
DRAM[14442] = 8'b10000110;
DRAM[14443] = 8'b10110100;
DRAM[14444] = 8'b11001011;
DRAM[14445] = 8'b11001000;
DRAM[14446] = 8'b11010011;
DRAM[14447] = 8'b11011010;
DRAM[14448] = 8'b11001110;
DRAM[14449] = 8'b10011110;
DRAM[14450] = 8'b01110110;
DRAM[14451] = 8'b01110010;
DRAM[14452] = 8'b01101001;
DRAM[14453] = 8'b01011110;
DRAM[14454] = 8'b01100010;
DRAM[14455] = 8'b01100010;
DRAM[14456] = 8'b01010000;
DRAM[14457] = 8'b01011110;
DRAM[14458] = 8'b01100111;
DRAM[14459] = 8'b01100100;
DRAM[14460] = 8'b01011111;
DRAM[14461] = 8'b01011111;
DRAM[14462] = 8'b01011101;
DRAM[14463] = 8'b01100010;
DRAM[14464] = 8'b00101000;
DRAM[14465] = 8'b00100110;
DRAM[14466] = 8'b01010010;
DRAM[14467] = 8'b10011011;
DRAM[14468] = 8'b10101010;
DRAM[14469] = 8'b10010111;
DRAM[14470] = 8'b01010010;
DRAM[14471] = 8'b01000001;
DRAM[14472] = 8'b10000100;
DRAM[14473] = 8'b10100010;
DRAM[14474] = 8'b10110000;
DRAM[14475] = 8'b10110001;
DRAM[14476] = 8'b10110001;
DRAM[14477] = 8'b10110000;
DRAM[14478] = 8'b10100011;
DRAM[14479] = 8'b10010101;
DRAM[14480] = 8'b10000101;
DRAM[14481] = 8'b01000001;
DRAM[14482] = 8'b00101010;
DRAM[14483] = 8'b00101000;
DRAM[14484] = 8'b00101110;
DRAM[14485] = 8'b01000101;
DRAM[14486] = 8'b01001000;
DRAM[14487] = 8'b00101110;
DRAM[14488] = 8'b00101110;
DRAM[14489] = 8'b00111110;
DRAM[14490] = 8'b00111010;
DRAM[14491] = 8'b00110011;
DRAM[14492] = 8'b00111010;
DRAM[14493] = 8'b00110101;
DRAM[14494] = 8'b00110111;
DRAM[14495] = 8'b00110010;
DRAM[14496] = 8'b00111010;
DRAM[14497] = 8'b01000100;
DRAM[14498] = 8'b00111110;
DRAM[14499] = 8'b01011000;
DRAM[14500] = 8'b00111101;
DRAM[14501] = 8'b10010000;
DRAM[14502] = 8'b01110001;
DRAM[14503] = 8'b01110011;
DRAM[14504] = 8'b01000101;
DRAM[14505] = 8'b01100010;
DRAM[14506] = 8'b01110011;
DRAM[14507] = 8'b01101100;
DRAM[14508] = 8'b01001011;
DRAM[14509] = 8'b00110110;
DRAM[14510] = 8'b00110010;
DRAM[14511] = 8'b00111011;
DRAM[14512] = 8'b00110101;
DRAM[14513] = 8'b00110010;
DRAM[14514] = 8'b00110011;
DRAM[14515] = 8'b00110000;
DRAM[14516] = 8'b01000110;
DRAM[14517] = 8'b01011010;
DRAM[14518] = 8'b01110000;
DRAM[14519] = 8'b01111100;
DRAM[14520] = 8'b10000000;
DRAM[14521] = 8'b01101011;
DRAM[14522] = 8'b01000000;
DRAM[14523] = 8'b01100110;
DRAM[14524] = 8'b10000001;
DRAM[14525] = 8'b10001001;
DRAM[14526] = 8'b10001100;
DRAM[14527] = 8'b10001011;
DRAM[14528] = 8'b10001110;
DRAM[14529] = 8'b10001011;
DRAM[14530] = 8'b10001010;
DRAM[14531] = 8'b10001000;
DRAM[14532] = 8'b10000111;
DRAM[14533] = 8'b10001011;
DRAM[14534] = 8'b10001000;
DRAM[14535] = 8'b10001010;
DRAM[14536] = 8'b10001110;
DRAM[14537] = 8'b10010010;
DRAM[14538] = 8'b10010011;
DRAM[14539] = 8'b10011001;
DRAM[14540] = 8'b10011001;
DRAM[14541] = 8'b10011110;
DRAM[14542] = 8'b10100100;
DRAM[14543] = 8'b10100101;
DRAM[14544] = 8'b10101100;
DRAM[14545] = 8'b10110100;
DRAM[14546] = 8'b10111011;
DRAM[14547] = 8'b11000010;
DRAM[14548] = 8'b11000110;
DRAM[14549] = 8'b11001011;
DRAM[14550] = 8'b11001111;
DRAM[14551] = 8'b11010001;
DRAM[14552] = 8'b11010100;
DRAM[14553] = 8'b11010100;
DRAM[14554] = 8'b11010110;
DRAM[14555] = 8'b10010100;
DRAM[14556] = 8'b10000110;
DRAM[14557] = 8'b10001010;
DRAM[14558] = 8'b10000111;
DRAM[14559] = 8'b10001011;
DRAM[14560] = 8'b10010000;
DRAM[14561] = 8'b10010010;
DRAM[14562] = 8'b10010010;
DRAM[14563] = 8'b10001111;
DRAM[14564] = 8'b10001110;
DRAM[14565] = 8'b10001101;
DRAM[14566] = 8'b10001000;
DRAM[14567] = 8'b10000110;
DRAM[14568] = 8'b10000111;
DRAM[14569] = 8'b10001000;
DRAM[14570] = 8'b10001001;
DRAM[14571] = 8'b10001111;
DRAM[14572] = 8'b10100100;
DRAM[14573] = 8'b10110110;
DRAM[14574] = 8'b11010100;
DRAM[14575] = 8'b11010111;
DRAM[14576] = 8'b11001000;
DRAM[14577] = 8'b10010001;
DRAM[14578] = 8'b01101110;
DRAM[14579] = 8'b01101011;
DRAM[14580] = 8'b01100000;
DRAM[14581] = 8'b01100000;
DRAM[14582] = 8'b01100100;
DRAM[14583] = 8'b01010100;
DRAM[14584] = 8'b01010010;
DRAM[14585] = 8'b01101001;
DRAM[14586] = 8'b01100100;
DRAM[14587] = 8'b01011111;
DRAM[14588] = 8'b01011000;
DRAM[14589] = 8'b01100010;
DRAM[14590] = 8'b01011111;
DRAM[14591] = 8'b01010110;
DRAM[14592] = 8'b00100100;
DRAM[14593] = 8'b00100110;
DRAM[14594] = 8'b01001010;
DRAM[14595] = 8'b10010110;
DRAM[14596] = 8'b10100111;
DRAM[14597] = 8'b10010111;
DRAM[14598] = 8'b01100000;
DRAM[14599] = 8'b01000011;
DRAM[14600] = 8'b01111110;
DRAM[14601] = 8'b10100000;
DRAM[14602] = 8'b10101111;
DRAM[14603] = 8'b10101110;
DRAM[14604] = 8'b10110001;
DRAM[14605] = 8'b10110010;
DRAM[14606] = 8'b10100101;
DRAM[14607] = 8'b10001110;
DRAM[14608] = 8'b10000111;
DRAM[14609] = 8'b01001011;
DRAM[14610] = 8'b00110100;
DRAM[14611] = 8'b00101110;
DRAM[14612] = 8'b01000000;
DRAM[14613] = 8'b00110110;
DRAM[14614] = 8'b00110001;
DRAM[14615] = 8'b00101111;
DRAM[14616] = 8'b00110011;
DRAM[14617] = 8'b01000000;
DRAM[14618] = 8'b00111100;
DRAM[14619] = 8'b01000010;
DRAM[14620] = 8'b00111101;
DRAM[14621] = 8'b00110101;
DRAM[14622] = 8'b00111101;
DRAM[14623] = 8'b00101110;
DRAM[14624] = 8'b00111101;
DRAM[14625] = 8'b01000001;
DRAM[14626] = 8'b00110000;
DRAM[14627] = 8'b01011100;
DRAM[14628] = 8'b01000011;
DRAM[14629] = 8'b00101111;
DRAM[14630] = 8'b01000111;
DRAM[14631] = 8'b01110000;
DRAM[14632] = 8'b00111100;
DRAM[14633] = 8'b01000011;
DRAM[14634] = 8'b01111100;
DRAM[14635] = 8'b10011010;
DRAM[14636] = 8'b00100111;
DRAM[14637] = 8'b00110001;
DRAM[14638] = 8'b00101100;
DRAM[14639] = 8'b00110110;
DRAM[14640] = 8'b00110001;
DRAM[14641] = 8'b00101100;
DRAM[14642] = 8'b00101111;
DRAM[14643] = 8'b00110101;
DRAM[14644] = 8'b01001011;
DRAM[14645] = 8'b01101010;
DRAM[14646] = 8'b01110101;
DRAM[14647] = 8'b01111110;
DRAM[14648] = 8'b01111011;
DRAM[14649] = 8'b01010000;
DRAM[14650] = 8'b01001101;
DRAM[14651] = 8'b01110010;
DRAM[14652] = 8'b10000100;
DRAM[14653] = 8'b10001001;
DRAM[14654] = 8'b10001010;
DRAM[14655] = 8'b10001110;
DRAM[14656] = 8'b10001111;
DRAM[14657] = 8'b10001111;
DRAM[14658] = 8'b10001100;
DRAM[14659] = 8'b10001110;
DRAM[14660] = 8'b10001001;
DRAM[14661] = 8'b10001000;
DRAM[14662] = 8'b10001011;
DRAM[14663] = 8'b10001100;
DRAM[14664] = 8'b10001110;
DRAM[14665] = 8'b10010001;
DRAM[14666] = 8'b10010011;
DRAM[14667] = 8'b10010111;
DRAM[14668] = 8'b10011000;
DRAM[14669] = 8'b10011011;
DRAM[14670] = 8'b10011110;
DRAM[14671] = 8'b10100101;
DRAM[14672] = 8'b10101100;
DRAM[14673] = 8'b10110010;
DRAM[14674] = 8'b10111000;
DRAM[14675] = 8'b11000000;
DRAM[14676] = 8'b11000110;
DRAM[14677] = 8'b11001001;
DRAM[14678] = 8'b11001111;
DRAM[14679] = 8'b11010010;
DRAM[14680] = 8'b11010011;
DRAM[14681] = 8'b11010101;
DRAM[14682] = 8'b11010100;
DRAM[14683] = 8'b11010100;
DRAM[14684] = 8'b10000101;
DRAM[14685] = 8'b01101110;
DRAM[14686] = 8'b01101100;
DRAM[14687] = 8'b01110010;
DRAM[14688] = 8'b01111010;
DRAM[14689] = 8'b10000100;
DRAM[14690] = 8'b10001011;
DRAM[14691] = 8'b10001111;
DRAM[14692] = 8'b10010001;
DRAM[14693] = 8'b10001111;
DRAM[14694] = 8'b10001100;
DRAM[14695] = 8'b10001001;
DRAM[14696] = 8'b10001110;
DRAM[14697] = 8'b10010101;
DRAM[14698] = 8'b10010001;
DRAM[14699] = 8'b10001010;
DRAM[14700] = 8'b10001010;
DRAM[14701] = 8'b10110101;
DRAM[14702] = 8'b11011000;
DRAM[14703] = 8'b11010110;
DRAM[14704] = 8'b10111100;
DRAM[14705] = 8'b10000000;
DRAM[14706] = 8'b01101111;
DRAM[14707] = 8'b01100010;
DRAM[14708] = 8'b01011100;
DRAM[14709] = 8'b01100010;
DRAM[14710] = 8'b01010110;
DRAM[14711] = 8'b01001111;
DRAM[14712] = 8'b01011111;
DRAM[14713] = 8'b01101000;
DRAM[14714] = 8'b01100001;
DRAM[14715] = 8'b01011011;
DRAM[14716] = 8'b01011101;
DRAM[14717] = 8'b01011110;
DRAM[14718] = 8'b01011111;
DRAM[14719] = 8'b01000110;
DRAM[14720] = 8'b00100010;
DRAM[14721] = 8'b00100100;
DRAM[14722] = 8'b01001001;
DRAM[14723] = 8'b10010001;
DRAM[14724] = 8'b10101010;
DRAM[14725] = 8'b10011110;
DRAM[14726] = 8'b01011100;
DRAM[14727] = 8'b01000110;
DRAM[14728] = 8'b01111100;
DRAM[14729] = 8'b10100010;
DRAM[14730] = 8'b10101100;
DRAM[14731] = 8'b10110000;
DRAM[14732] = 8'b10110010;
DRAM[14733] = 8'b10110001;
DRAM[14734] = 8'b10100110;
DRAM[14735] = 8'b10001100;
DRAM[14736] = 8'b01110110;
DRAM[14737] = 8'b01001011;
DRAM[14738] = 8'b00111000;
DRAM[14739] = 8'b00101110;
DRAM[14740] = 8'b00110111;
DRAM[14741] = 8'b00110100;
DRAM[14742] = 8'b00110000;
DRAM[14743] = 8'b00110000;
DRAM[14744] = 8'b00111100;
DRAM[14745] = 8'b00111111;
DRAM[14746] = 8'b00110110;
DRAM[14747] = 8'b01001010;
DRAM[14748] = 8'b00110100;
DRAM[14749] = 8'b00101110;
DRAM[14750] = 8'b00110010;
DRAM[14751] = 8'b00101000;
DRAM[14752] = 8'b01000000;
DRAM[14753] = 8'b00110011;
DRAM[14754] = 8'b00111000;
DRAM[14755] = 8'b01101000;
DRAM[14756] = 8'b01101000;
DRAM[14757] = 8'b00111101;
DRAM[14758] = 8'b00110001;
DRAM[14759] = 8'b01001111;
DRAM[14760] = 8'b01001000;
DRAM[14761] = 8'b01011010;
DRAM[14762] = 8'b01011101;
DRAM[14763] = 8'b01100100;
DRAM[14764] = 8'b00101100;
DRAM[14765] = 8'b00110101;
DRAM[14766] = 8'b00101111;
DRAM[14767] = 8'b00110000;
DRAM[14768] = 8'b00110000;
DRAM[14769] = 8'b00101000;
DRAM[14770] = 8'b00110001;
DRAM[14771] = 8'b01000010;
DRAM[14772] = 8'b01010111;
DRAM[14773] = 8'b01110000;
DRAM[14774] = 8'b01110111;
DRAM[14775] = 8'b01111100;
DRAM[14776] = 8'b01110011;
DRAM[14777] = 8'b00110110;
DRAM[14778] = 8'b01011010;
DRAM[14779] = 8'b10000100;
DRAM[14780] = 8'b10000110;
DRAM[14781] = 8'b10001000;
DRAM[14782] = 8'b10001011;
DRAM[14783] = 8'b10001111;
DRAM[14784] = 8'b10010000;
DRAM[14785] = 8'b10001111;
DRAM[14786] = 8'b10001101;
DRAM[14787] = 8'b10001111;
DRAM[14788] = 8'b10001011;
DRAM[14789] = 8'b10000111;
DRAM[14790] = 8'b10001010;
DRAM[14791] = 8'b10001011;
DRAM[14792] = 8'b10001110;
DRAM[14793] = 8'b10010001;
DRAM[14794] = 8'b10010100;
DRAM[14795] = 8'b10010110;
DRAM[14796] = 8'b10011000;
DRAM[14797] = 8'b10011001;
DRAM[14798] = 8'b10100010;
DRAM[14799] = 8'b10100011;
DRAM[14800] = 8'b10101001;
DRAM[14801] = 8'b10101011;
DRAM[14802] = 8'b10110110;
DRAM[14803] = 8'b10111101;
DRAM[14804] = 8'b11000010;
DRAM[14805] = 8'b11001001;
DRAM[14806] = 8'b11001110;
DRAM[14807] = 8'b11010001;
DRAM[14808] = 8'b11010011;
DRAM[14809] = 8'b11010100;
DRAM[14810] = 8'b11010111;
DRAM[14811] = 8'b11011010;
DRAM[14812] = 8'b10001101;
DRAM[14813] = 8'b01010000;
DRAM[14814] = 8'b01010000;
DRAM[14815] = 8'b01010000;
DRAM[14816] = 8'b01011010;
DRAM[14817] = 8'b01100111;
DRAM[14818] = 8'b01110000;
DRAM[14819] = 8'b01111010;
DRAM[14820] = 8'b01111111;
DRAM[14821] = 8'b10000101;
DRAM[14822] = 8'b10001000;
DRAM[14823] = 8'b10001111;
DRAM[14824] = 8'b10010101;
DRAM[14825] = 8'b10011010;
DRAM[14826] = 8'b10001101;
DRAM[14827] = 8'b10000011;
DRAM[14828] = 8'b10010000;
DRAM[14829] = 8'b11000110;
DRAM[14830] = 8'b11011011;
DRAM[14831] = 8'b11010000;
DRAM[14832] = 8'b10100110;
DRAM[14833] = 8'b01110101;
DRAM[14834] = 8'b01100010;
DRAM[14835] = 8'b01010101;
DRAM[14836] = 8'b01011100;
DRAM[14837] = 8'b01011101;
DRAM[14838] = 8'b01001000;
DRAM[14839] = 8'b01010111;
DRAM[14840] = 8'b01101001;
DRAM[14841] = 8'b01100001;
DRAM[14842] = 8'b01011110;
DRAM[14843] = 8'b01011010;
DRAM[14844] = 8'b01101000;
DRAM[14845] = 8'b01011100;
DRAM[14846] = 8'b01010100;
DRAM[14847] = 8'b00111011;
DRAM[14848] = 8'b00100010;
DRAM[14849] = 8'b00100001;
DRAM[14850] = 8'b00111000;
DRAM[14851] = 8'b10011000;
DRAM[14852] = 8'b10101110;
DRAM[14853] = 8'b10100101;
DRAM[14854] = 8'b01101101;
DRAM[14855] = 8'b01000000;
DRAM[14856] = 8'b01111001;
DRAM[14857] = 8'b10011101;
DRAM[14858] = 8'b10101100;
DRAM[14859] = 8'b10101111;
DRAM[14860] = 8'b10110000;
DRAM[14861] = 8'b10110011;
DRAM[14862] = 8'b10101000;
DRAM[14863] = 8'b10010010;
DRAM[14864] = 8'b01110011;
DRAM[14865] = 8'b01010001;
DRAM[14866] = 8'b00110010;
DRAM[14867] = 8'b00110001;
DRAM[14868] = 8'b00101101;
DRAM[14869] = 8'b00101100;
DRAM[14870] = 8'b00101101;
DRAM[14871] = 8'b00111111;
DRAM[14872] = 8'b00101110;
DRAM[14873] = 8'b00111011;
DRAM[14874] = 8'b00110011;
DRAM[14875] = 8'b01000100;
DRAM[14876] = 8'b00110111;
DRAM[14877] = 8'b00101110;
DRAM[14878] = 8'b00101101;
DRAM[14879] = 8'b00110011;
DRAM[14880] = 8'b00110011;
DRAM[14881] = 8'b00110110;
DRAM[14882] = 8'b01010001;
DRAM[14883] = 8'b01011110;
DRAM[14884] = 8'b10000100;
DRAM[14885] = 8'b01010110;
DRAM[14886] = 8'b00111110;
DRAM[14887] = 8'b01000100;
DRAM[14888] = 8'b01000110;
DRAM[14889] = 8'b01101110;
DRAM[14890] = 8'b01000000;
DRAM[14891] = 8'b01001010;
DRAM[14892] = 8'b00110010;
DRAM[14893] = 8'b00101010;
DRAM[14894] = 8'b00110011;
DRAM[14895] = 8'b00101100;
DRAM[14896] = 8'b00101100;
DRAM[14897] = 8'b00101001;
DRAM[14898] = 8'b00111001;
DRAM[14899] = 8'b01001111;
DRAM[14900] = 8'b01101001;
DRAM[14901] = 8'b01110110;
DRAM[14902] = 8'b01110101;
DRAM[14903] = 8'b01110110;
DRAM[14904] = 8'b01010100;
DRAM[14905] = 8'b01000000;
DRAM[14906] = 8'b01101100;
DRAM[14907] = 8'b10000101;
DRAM[14908] = 8'b10000111;
DRAM[14909] = 8'b10000111;
DRAM[14910] = 8'b10001100;
DRAM[14911] = 8'b10001110;
DRAM[14912] = 8'b10010001;
DRAM[14913] = 8'b10001011;
DRAM[14914] = 8'b10001110;
DRAM[14915] = 8'b10001011;
DRAM[14916] = 8'b10001100;
DRAM[14917] = 8'b10001010;
DRAM[14918] = 8'b10000110;
DRAM[14919] = 8'b10001001;
DRAM[14920] = 8'b10001010;
DRAM[14921] = 8'b10010000;
DRAM[14922] = 8'b10010001;
DRAM[14923] = 8'b10010100;
DRAM[14924] = 8'b10010101;
DRAM[14925] = 8'b10011011;
DRAM[14926] = 8'b10011110;
DRAM[14927] = 8'b10100010;
DRAM[14928] = 8'b10101000;
DRAM[14929] = 8'b10101010;
DRAM[14930] = 8'b10110001;
DRAM[14931] = 8'b10111011;
DRAM[14932] = 8'b11000001;
DRAM[14933] = 8'b11001000;
DRAM[14934] = 8'b11001100;
DRAM[14935] = 8'b11001111;
DRAM[14936] = 8'b11010100;
DRAM[14937] = 8'b11010110;
DRAM[14938] = 8'b11010111;
DRAM[14939] = 8'b11011010;
DRAM[14940] = 8'b10010011;
DRAM[14941] = 8'b01010011;
DRAM[14942] = 8'b01010100;
DRAM[14943] = 8'b01001100;
DRAM[14944] = 8'b01001010;
DRAM[14945] = 8'b01001110;
DRAM[14946] = 8'b01010001;
DRAM[14947] = 8'b01010100;
DRAM[14948] = 8'b01011001;
DRAM[14949] = 8'b01100011;
DRAM[14950] = 8'b01101010;
DRAM[14951] = 8'b01111100;
DRAM[14952] = 8'b10010001;
DRAM[14953] = 8'b10011110;
DRAM[14954] = 8'b10010001;
DRAM[14955] = 8'b10001101;
DRAM[14956] = 8'b10011001;
DRAM[14957] = 8'b11010001;
DRAM[14958] = 8'b11011011;
DRAM[14959] = 8'b11000011;
DRAM[14960] = 8'b10001011;
DRAM[14961] = 8'b01100001;
DRAM[14962] = 8'b01001111;
DRAM[14963] = 8'b01001110;
DRAM[14964] = 8'b01011011;
DRAM[14965] = 8'b01010010;
DRAM[14966] = 8'b01010010;
DRAM[14967] = 8'b01100111;
DRAM[14968] = 8'b01100010;
DRAM[14969] = 8'b01011100;
DRAM[14970] = 8'b01011100;
DRAM[14971] = 8'b01100001;
DRAM[14972] = 8'b01100111;
DRAM[14973] = 8'b01011110;
DRAM[14974] = 8'b01000011;
DRAM[14975] = 8'b00110100;
DRAM[14976] = 8'b00100110;
DRAM[14977] = 8'b00100101;
DRAM[14978] = 8'b00110110;
DRAM[14979] = 8'b10010110;
DRAM[14980] = 8'b10101111;
DRAM[14981] = 8'b10101000;
DRAM[14982] = 8'b10000000;
DRAM[14983] = 8'b01000010;
DRAM[14984] = 8'b01110110;
DRAM[14985] = 8'b10011110;
DRAM[14986] = 8'b10101011;
DRAM[14987] = 8'b10110000;
DRAM[14988] = 8'b10110000;
DRAM[14989] = 8'b10110100;
DRAM[14990] = 8'b10101010;
DRAM[14991] = 8'b10000110;
DRAM[14992] = 8'b01101010;
DRAM[14993] = 8'b01010100;
DRAM[14994] = 8'b00101111;
DRAM[14995] = 8'b00110010;
DRAM[14996] = 8'b00101011;
DRAM[14997] = 8'b00101010;
DRAM[14998] = 8'b01000001;
DRAM[14999] = 8'b00111010;
DRAM[15000] = 8'b00101111;
DRAM[15001] = 8'b00111100;
DRAM[15002] = 8'b00110100;
DRAM[15003] = 8'b00111111;
DRAM[15004] = 8'b00111111;
DRAM[15005] = 8'b00111011;
DRAM[15006] = 8'b00110000;
DRAM[15007] = 8'b00110100;
DRAM[15008] = 8'b00111010;
DRAM[15009] = 8'b00101010;
DRAM[15010] = 8'b00101101;
DRAM[15011] = 8'b01010000;
DRAM[15012] = 8'b01110000;
DRAM[15013] = 8'b10001000;
DRAM[15014] = 8'b01101110;
DRAM[15015] = 8'b01101000;
DRAM[15016] = 8'b01101010;
DRAM[15017] = 8'b00111001;
DRAM[15018] = 8'b00101110;
DRAM[15019] = 8'b00110011;
DRAM[15020] = 8'b00110111;
DRAM[15021] = 8'b00101111;
DRAM[15022] = 8'b00101011;
DRAM[15023] = 8'b00101000;
DRAM[15024] = 8'b00101000;
DRAM[15025] = 8'b00110000;
DRAM[15026] = 8'b01000100;
DRAM[15027] = 8'b01011100;
DRAM[15028] = 8'b01101110;
DRAM[15029] = 8'b01110101;
DRAM[15030] = 8'b01111000;
DRAM[15031] = 8'b01101000;
DRAM[15032] = 8'b00101011;
DRAM[15033] = 8'b01011101;
DRAM[15034] = 8'b10000000;
DRAM[15035] = 8'b10000111;
DRAM[15036] = 8'b10000110;
DRAM[15037] = 8'b10001010;
DRAM[15038] = 8'b10001011;
DRAM[15039] = 8'b10001101;
DRAM[15040] = 8'b10001110;
DRAM[15041] = 8'b10001101;
DRAM[15042] = 8'b10001111;
DRAM[15043] = 8'b10001100;
DRAM[15044] = 8'b10001010;
DRAM[15045] = 8'b10001001;
DRAM[15046] = 8'b10000111;
DRAM[15047] = 8'b10000111;
DRAM[15048] = 8'b10001001;
DRAM[15049] = 8'b10001011;
DRAM[15050] = 8'b10010001;
DRAM[15051] = 8'b10010011;
DRAM[15052] = 8'b10010111;
DRAM[15053] = 8'b10010110;
DRAM[15054] = 8'b10011100;
DRAM[15055] = 8'b10011100;
DRAM[15056] = 8'b10100101;
DRAM[15057] = 8'b10101001;
DRAM[15058] = 8'b10110001;
DRAM[15059] = 8'b10111000;
DRAM[15060] = 8'b10111110;
DRAM[15061] = 8'b11000110;
DRAM[15062] = 8'b11001010;
DRAM[15063] = 8'b11001111;
DRAM[15064] = 8'b11010001;
DRAM[15065] = 8'b11010100;
DRAM[15066] = 8'b11010101;
DRAM[15067] = 8'b11011010;
DRAM[15068] = 8'b11000011;
DRAM[15069] = 8'b01010000;
DRAM[15070] = 8'b01100011;
DRAM[15071] = 8'b01100000;
DRAM[15072] = 8'b01011000;
DRAM[15073] = 8'b01010011;
DRAM[15074] = 8'b01001010;
DRAM[15075] = 8'b01000010;
DRAM[15076] = 8'b00111010;
DRAM[15077] = 8'b00111001;
DRAM[15078] = 8'b00111001;
DRAM[15079] = 8'b01001010;
DRAM[15080] = 8'b01101000;
DRAM[15081] = 8'b10001111;
DRAM[15082] = 8'b10110110;
DRAM[15083] = 8'b10100001;
DRAM[15084] = 8'b10110001;
DRAM[15085] = 8'b11010110;
DRAM[15086] = 8'b11010101;
DRAM[15087] = 8'b10101010;
DRAM[15088] = 8'b01101101;
DRAM[15089] = 8'b01001001;
DRAM[15090] = 8'b00111011;
DRAM[15091] = 8'b01010000;
DRAM[15092] = 8'b01010000;
DRAM[15093] = 8'b01010101;
DRAM[15094] = 8'b01100100;
DRAM[15095] = 8'b01100100;
DRAM[15096] = 8'b01011001;
DRAM[15097] = 8'b01011010;
DRAM[15098] = 8'b01011010;
DRAM[15099] = 8'b01100101;
DRAM[15100] = 8'b01100010;
DRAM[15101] = 8'b01010111;
DRAM[15102] = 8'b00111100;
DRAM[15103] = 8'b00110111;
DRAM[15104] = 8'b00111010;
DRAM[15105] = 8'b01000001;
DRAM[15106] = 8'b01000111;
DRAM[15107] = 8'b10001110;
DRAM[15108] = 8'b10110011;
DRAM[15109] = 8'b10110010;
DRAM[15110] = 8'b10000110;
DRAM[15111] = 8'b01000101;
DRAM[15112] = 8'b01110101;
DRAM[15113] = 8'b10011100;
DRAM[15114] = 8'b10101101;
DRAM[15115] = 8'b10110000;
DRAM[15116] = 8'b10101110;
DRAM[15117] = 8'b10110110;
DRAM[15118] = 8'b10101010;
DRAM[15119] = 8'b01111010;
DRAM[15120] = 8'b01110000;
DRAM[15121] = 8'b00111110;
DRAM[15122] = 8'b00101110;
DRAM[15123] = 8'b00110011;
DRAM[15124] = 8'b00110100;
DRAM[15125] = 8'b00111000;
DRAM[15126] = 8'b00110100;
DRAM[15127] = 8'b00111000;
DRAM[15128] = 8'b00101110;
DRAM[15129] = 8'b00111010;
DRAM[15130] = 8'b00111000;
DRAM[15131] = 8'b00111111;
DRAM[15132] = 8'b00111011;
DRAM[15133] = 8'b00110100;
DRAM[15134] = 8'b00110110;
DRAM[15135] = 8'b00101101;
DRAM[15136] = 8'b00101110;
DRAM[15137] = 8'b00111000;
DRAM[15138] = 8'b00110100;
DRAM[15139] = 8'b00101010;
DRAM[15140] = 8'b01010010;
DRAM[15141] = 8'b10010100;
DRAM[15142] = 8'b10000001;
DRAM[15143] = 8'b01100000;
DRAM[15144] = 8'b01100000;
DRAM[15145] = 8'b01100011;
DRAM[15146] = 8'b00101000;
DRAM[15147] = 8'b00110001;
DRAM[15148] = 8'b00101010;
DRAM[15149] = 8'b00101111;
DRAM[15150] = 8'b00110000;
DRAM[15151] = 8'b00101010;
DRAM[15152] = 8'b00101100;
DRAM[15153] = 8'b00111000;
DRAM[15154] = 8'b01001111;
DRAM[15155] = 8'b01100110;
DRAM[15156] = 8'b01110001;
DRAM[15157] = 8'b01110110;
DRAM[15158] = 8'b01110011;
DRAM[15159] = 8'b00110011;
DRAM[15160] = 8'b01000000;
DRAM[15161] = 8'b01110111;
DRAM[15162] = 8'b10000011;
DRAM[15163] = 8'b10001001;
DRAM[15164] = 8'b10001001;
DRAM[15165] = 8'b10001010;
DRAM[15166] = 8'b10001010;
DRAM[15167] = 8'b10001011;
DRAM[15168] = 8'b10001010;
DRAM[15169] = 8'b10010001;
DRAM[15170] = 8'b10010000;
DRAM[15171] = 8'b10001110;
DRAM[15172] = 8'b10001100;
DRAM[15173] = 8'b10001100;
DRAM[15174] = 8'b10001011;
DRAM[15175] = 8'b10001000;
DRAM[15176] = 8'b10001011;
DRAM[15177] = 8'b10001010;
DRAM[15178] = 8'b10001100;
DRAM[15179] = 8'b10001111;
DRAM[15180] = 8'b10010100;
DRAM[15181] = 8'b10010111;
DRAM[15182] = 8'b10011011;
DRAM[15183] = 8'b10011110;
DRAM[15184] = 8'b10100000;
DRAM[15185] = 8'b10100111;
DRAM[15186] = 8'b10110001;
DRAM[15187] = 8'b10110100;
DRAM[15188] = 8'b10111011;
DRAM[15189] = 8'b11000011;
DRAM[15190] = 8'b11001000;
DRAM[15191] = 8'b11001101;
DRAM[15192] = 8'b11010000;
DRAM[15193] = 8'b11010011;
DRAM[15194] = 8'b11010100;
DRAM[15195] = 8'b11011000;
DRAM[15196] = 8'b11011001;
DRAM[15197] = 8'b01011100;
DRAM[15198] = 8'b01100001;
DRAM[15199] = 8'b01101001;
DRAM[15200] = 8'b01100110;
DRAM[15201] = 8'b01011101;
DRAM[15202] = 8'b01011000;
DRAM[15203] = 8'b01001100;
DRAM[15204] = 8'b00111111;
DRAM[15205] = 8'b00110010;
DRAM[15206] = 8'b00101000;
DRAM[15207] = 8'b00101001;
DRAM[15208] = 8'b01001110;
DRAM[15209] = 8'b10111000;
DRAM[15210] = 8'b11000111;
DRAM[15211] = 8'b10100011;
DRAM[15212] = 8'b10111100;
DRAM[15213] = 8'b11010110;
DRAM[15214] = 8'b11001011;
DRAM[15215] = 8'b10000111;
DRAM[15216] = 8'b01000110;
DRAM[15217] = 8'b00111100;
DRAM[15218] = 8'b01001010;
DRAM[15219] = 8'b01001110;
DRAM[15220] = 8'b01000111;
DRAM[15221] = 8'b01011110;
DRAM[15222] = 8'b01101000;
DRAM[15223] = 8'b01011100;
DRAM[15224] = 8'b01010111;
DRAM[15225] = 8'b01010100;
DRAM[15226] = 8'b01011110;
DRAM[15227] = 8'b01101010;
DRAM[15228] = 8'b01100000;
DRAM[15229] = 8'b01001010;
DRAM[15230] = 8'b00111101;
DRAM[15231] = 8'b00110110;
DRAM[15232] = 8'b01011011;
DRAM[15233] = 8'b01011000;
DRAM[15234] = 8'b01100000;
DRAM[15235] = 8'b10001010;
DRAM[15236] = 8'b10110000;
DRAM[15237] = 8'b10110011;
DRAM[15238] = 8'b10001101;
DRAM[15239] = 8'b01001110;
DRAM[15240] = 8'b01110110;
DRAM[15241] = 8'b10011100;
DRAM[15242] = 8'b10101101;
DRAM[15243] = 8'b10110001;
DRAM[15244] = 8'b10101110;
DRAM[15245] = 8'b10110110;
DRAM[15246] = 8'b10101010;
DRAM[15247] = 8'b01111100;
DRAM[15248] = 8'b01111000;
DRAM[15249] = 8'b01001000;
DRAM[15250] = 8'b00101100;
DRAM[15251] = 8'b00110101;
DRAM[15252] = 8'b00111011;
DRAM[15253] = 8'b00110010;
DRAM[15254] = 8'b00110000;
DRAM[15255] = 8'b00110011;
DRAM[15256] = 8'b00110000;
DRAM[15257] = 8'b00110011;
DRAM[15258] = 8'b00111111;
DRAM[15259] = 8'b00111010;
DRAM[15260] = 8'b00111100;
DRAM[15261] = 8'b00111110;
DRAM[15262] = 8'b00101111;
DRAM[15263] = 8'b00101011;
DRAM[15264] = 8'b00110010;
DRAM[15265] = 8'b00110100;
DRAM[15266] = 8'b01000010;
DRAM[15267] = 8'b00110011;
DRAM[15268] = 8'b00101101;
DRAM[15269] = 8'b01010010;
DRAM[15270] = 8'b10001011;
DRAM[15271] = 8'b10001010;
DRAM[15272] = 8'b01011100;
DRAM[15273] = 8'b01110000;
DRAM[15274] = 8'b00110000;
DRAM[15275] = 8'b00101110;
DRAM[15276] = 8'b00101010;
DRAM[15277] = 8'b00101000;
DRAM[15278] = 8'b00100111;
DRAM[15279] = 8'b00101101;
DRAM[15280] = 8'b00101111;
DRAM[15281] = 8'b01001011;
DRAM[15282] = 8'b01011010;
DRAM[15283] = 8'b01110011;
DRAM[15284] = 8'b01111000;
DRAM[15285] = 8'b01110100;
DRAM[15286] = 8'b00110101;
DRAM[15287] = 8'b00110010;
DRAM[15288] = 8'b01100110;
DRAM[15289] = 8'b10000000;
DRAM[15290] = 8'b10000010;
DRAM[15291] = 8'b10000101;
DRAM[15292] = 8'b10001000;
DRAM[15293] = 8'b10001011;
DRAM[15294] = 8'b10001100;
DRAM[15295] = 8'b10001100;
DRAM[15296] = 8'b10001100;
DRAM[15297] = 8'b10001110;
DRAM[15298] = 8'b10001111;
DRAM[15299] = 8'b10001111;
DRAM[15300] = 8'b10001111;
DRAM[15301] = 8'b10001100;
DRAM[15302] = 8'b10001001;
DRAM[15303] = 8'b10001001;
DRAM[15304] = 8'b10001001;
DRAM[15305] = 8'b10001100;
DRAM[15306] = 8'b10001000;
DRAM[15307] = 8'b10001101;
DRAM[15308] = 8'b10010001;
DRAM[15309] = 8'b10010011;
DRAM[15310] = 8'b10011000;
DRAM[15311] = 8'b10011010;
DRAM[15312] = 8'b10100000;
DRAM[15313] = 8'b10100110;
DRAM[15314] = 8'b10101010;
DRAM[15315] = 8'b10110000;
DRAM[15316] = 8'b10111001;
DRAM[15317] = 8'b11000000;
DRAM[15318] = 8'b11000110;
DRAM[15319] = 8'b11001011;
DRAM[15320] = 8'b11001110;
DRAM[15321] = 8'b11010000;
DRAM[15322] = 8'b11010100;
DRAM[15323] = 8'b11010111;
DRAM[15324] = 8'b11011000;
DRAM[15325] = 8'b10000110;
DRAM[15326] = 8'b01011110;
DRAM[15327] = 8'b01101000;
DRAM[15328] = 8'b01101010;
DRAM[15329] = 8'b01100100;
DRAM[15330] = 8'b01011110;
DRAM[15331] = 8'b01011001;
DRAM[15332] = 8'b01001110;
DRAM[15333] = 8'b01000000;
DRAM[15334] = 8'b00110000;
DRAM[15335] = 8'b00101000;
DRAM[15336] = 8'b01001011;
DRAM[15337] = 8'b10111111;
DRAM[15338] = 8'b11000111;
DRAM[15339] = 8'b10100101;
DRAM[15340] = 8'b11000110;
DRAM[15341] = 8'b11001100;
DRAM[15342] = 8'b10100110;
DRAM[15343] = 8'b01001010;
DRAM[15344] = 8'b00111000;
DRAM[15345] = 8'b01000000;
DRAM[15346] = 8'b01001010;
DRAM[15347] = 8'b01000111;
DRAM[15348] = 8'b01010110;
DRAM[15349] = 8'b01101011;
DRAM[15350] = 8'b01011101;
DRAM[15351] = 8'b01010001;
DRAM[15352] = 8'b01010000;
DRAM[15353] = 8'b01010110;
DRAM[15354] = 8'b01100111;
DRAM[15355] = 8'b01101101;
DRAM[15356] = 8'b01011100;
DRAM[15357] = 8'b01010001;
DRAM[15358] = 8'b00111111;
DRAM[15359] = 8'b00111100;
DRAM[15360] = 8'b01011000;
DRAM[15361] = 8'b01100000;
DRAM[15362] = 8'b01101111;
DRAM[15363] = 8'b10010001;
DRAM[15364] = 8'b10110000;
DRAM[15365] = 8'b10110101;
DRAM[15366] = 8'b10010111;
DRAM[15367] = 8'b01010111;
DRAM[15368] = 8'b01110011;
DRAM[15369] = 8'b10011101;
DRAM[15370] = 8'b10101101;
DRAM[15371] = 8'b10110010;
DRAM[15372] = 8'b10110010;
DRAM[15373] = 8'b10110111;
DRAM[15374] = 8'b10101110;
DRAM[15375] = 8'b01110111;
DRAM[15376] = 8'b01110110;
DRAM[15377] = 8'b01000010;
DRAM[15378] = 8'b00101111;
DRAM[15379] = 8'b00110000;
DRAM[15380] = 8'b00110001;
DRAM[15381] = 8'b00101111;
DRAM[15382] = 8'b00101110;
DRAM[15383] = 8'b00111001;
DRAM[15384] = 8'b00110100;
DRAM[15385] = 8'b00110001;
DRAM[15386] = 8'b00101110;
DRAM[15387] = 8'b01000010;
DRAM[15388] = 8'b00110110;
DRAM[15389] = 8'b00111101;
DRAM[15390] = 8'b00111011;
DRAM[15391] = 8'b00101101;
DRAM[15392] = 8'b00110110;
DRAM[15393] = 8'b00111110;
DRAM[15394] = 8'b00111011;
DRAM[15395] = 8'b00111001;
DRAM[15396] = 8'b01001001;
DRAM[15397] = 8'b01000001;
DRAM[15398] = 8'b01010010;
DRAM[15399] = 8'b01011010;
DRAM[15400] = 8'b10001000;
DRAM[15401] = 8'b00110001;
DRAM[15402] = 8'b00101110;
DRAM[15403] = 8'b00110000;
DRAM[15404] = 8'b00101110;
DRAM[15405] = 8'b00101011;
DRAM[15406] = 8'b00100111;
DRAM[15407] = 8'b00101111;
DRAM[15408] = 8'b01000000;
DRAM[15409] = 8'b01010100;
DRAM[15410] = 8'b01100101;
DRAM[15411] = 8'b01110110;
DRAM[15412] = 8'b01101100;
DRAM[15413] = 8'b00110111;
DRAM[15414] = 8'b00110011;
DRAM[15415] = 8'b01100100;
DRAM[15416] = 8'b01111011;
DRAM[15417] = 8'b10000001;
DRAM[15418] = 8'b10000011;
DRAM[15419] = 8'b10000110;
DRAM[15420] = 8'b10001001;
DRAM[15421] = 8'b10001100;
DRAM[15422] = 8'b10001010;
DRAM[15423] = 8'b10001011;
DRAM[15424] = 8'b10001011;
DRAM[15425] = 8'b10001110;
DRAM[15426] = 8'b10001111;
DRAM[15427] = 8'b10001011;
DRAM[15428] = 8'b10001111;
DRAM[15429] = 8'b10001110;
DRAM[15430] = 8'b10001111;
DRAM[15431] = 8'b10001000;
DRAM[15432] = 8'b10001011;
DRAM[15433] = 8'b10001011;
DRAM[15434] = 8'b10001101;
DRAM[15435] = 8'b10001101;
DRAM[15436] = 8'b10010001;
DRAM[15437] = 8'b10010011;
DRAM[15438] = 8'b10010101;
DRAM[15439] = 8'b10011001;
DRAM[15440] = 8'b10100000;
DRAM[15441] = 8'b10100100;
DRAM[15442] = 8'b10100100;
DRAM[15443] = 8'b10101101;
DRAM[15444] = 8'b10110110;
DRAM[15445] = 8'b10111101;
DRAM[15446] = 8'b11000010;
DRAM[15447] = 8'b11001001;
DRAM[15448] = 8'b11001110;
DRAM[15449] = 8'b11010000;
DRAM[15450] = 8'b11010010;
DRAM[15451] = 8'b11010011;
DRAM[15452] = 8'b11010111;
DRAM[15453] = 8'b10101011;
DRAM[15454] = 8'b01010101;
DRAM[15455] = 8'b01100111;
DRAM[15456] = 8'b01101011;
DRAM[15457] = 8'b01101000;
DRAM[15458] = 8'b01100100;
DRAM[15459] = 8'b01100000;
DRAM[15460] = 8'b01010101;
DRAM[15461] = 8'b01001011;
DRAM[15462] = 8'b01000001;
DRAM[15463] = 8'b00111101;
DRAM[15464] = 8'b01010000;
DRAM[15465] = 8'b10110010;
DRAM[15466] = 8'b11001011;
DRAM[15467] = 8'b11000100;
DRAM[15468] = 8'b10110111;
DRAM[15469] = 8'b10011100;
DRAM[15470] = 8'b01010010;
DRAM[15471] = 8'b00110100;
DRAM[15472] = 8'b00111000;
DRAM[15473] = 8'b01000100;
DRAM[15474] = 8'b01000001;
DRAM[15475] = 8'b01010101;
DRAM[15476] = 8'b01100111;
DRAM[15477] = 8'b01100011;
DRAM[15478] = 8'b01001110;
DRAM[15479] = 8'b01001111;
DRAM[15480] = 8'b01010000;
DRAM[15481] = 8'b01100010;
DRAM[15482] = 8'b01110000;
DRAM[15483] = 8'b01100100;
DRAM[15484] = 8'b01011010;
DRAM[15485] = 8'b01001010;
DRAM[15486] = 8'b00111011;
DRAM[15487] = 8'b01000011;
DRAM[15488] = 8'b01001010;
DRAM[15489] = 8'b01101011;
DRAM[15490] = 8'b01110011;
DRAM[15491] = 8'b10001010;
DRAM[15492] = 8'b10101100;
DRAM[15493] = 8'b10110000;
DRAM[15494] = 8'b10010100;
DRAM[15495] = 8'b01011101;
DRAM[15496] = 8'b01110101;
DRAM[15497] = 8'b10011011;
DRAM[15498] = 8'b10101010;
DRAM[15499] = 8'b10110001;
DRAM[15500] = 8'b10110011;
DRAM[15501] = 8'b10110110;
DRAM[15502] = 8'b10101011;
DRAM[15503] = 8'b01110010;
DRAM[15504] = 8'b01110100;
DRAM[15505] = 8'b00111100;
DRAM[15506] = 8'b00101100;
DRAM[15507] = 8'b00110011;
DRAM[15508] = 8'b00110111;
DRAM[15509] = 8'b00110110;
DRAM[15510] = 8'b00110101;
DRAM[15511] = 8'b00111010;
DRAM[15512] = 8'b00110000;
DRAM[15513] = 8'b00101010;
DRAM[15514] = 8'b00111000;
DRAM[15515] = 8'b01011001;
DRAM[15516] = 8'b00110011;
DRAM[15517] = 8'b01001100;
DRAM[15518] = 8'b01001000;
DRAM[15519] = 8'b00101100;
DRAM[15520] = 8'b00111100;
DRAM[15521] = 8'b01001100;
DRAM[15522] = 8'b00111010;
DRAM[15523] = 8'b01001000;
DRAM[15524] = 8'b01000100;
DRAM[15525] = 8'b01000101;
DRAM[15526] = 8'b01100000;
DRAM[15527] = 8'b01100001;
DRAM[15528] = 8'b00111010;
DRAM[15529] = 8'b01000110;
DRAM[15530] = 8'b00101010;
DRAM[15531] = 8'b00101101;
DRAM[15532] = 8'b00101100;
DRAM[15533] = 8'b00100100;
DRAM[15534] = 8'b00100111;
DRAM[15535] = 8'b00110101;
DRAM[15536] = 8'b01001101;
DRAM[15537] = 8'b01011111;
DRAM[15538] = 8'b01011011;
DRAM[15539] = 8'b01000111;
DRAM[15540] = 8'b00101111;
DRAM[15541] = 8'b01000111;
DRAM[15542] = 8'b01101000;
DRAM[15543] = 8'b01110100;
DRAM[15544] = 8'b01111111;
DRAM[15545] = 8'b10000011;
DRAM[15546] = 8'b10000100;
DRAM[15547] = 8'b10001010;
DRAM[15548] = 8'b10001000;
DRAM[15549] = 8'b10001011;
DRAM[15550] = 8'b10001010;
DRAM[15551] = 8'b10001101;
DRAM[15552] = 8'b10001100;
DRAM[15553] = 8'b10001110;
DRAM[15554] = 8'b10001110;
DRAM[15555] = 8'b10001101;
DRAM[15556] = 8'b10001111;
DRAM[15557] = 8'b10001110;
DRAM[15558] = 8'b10001111;
DRAM[15559] = 8'b10001100;
DRAM[15560] = 8'b10001101;
DRAM[15561] = 8'b10001100;
DRAM[15562] = 8'b10001011;
DRAM[15563] = 8'b10001100;
DRAM[15564] = 8'b10001111;
DRAM[15565] = 8'b10010011;
DRAM[15566] = 8'b10010011;
DRAM[15567] = 8'b10011010;
DRAM[15568] = 8'b10011100;
DRAM[15569] = 8'b10100000;
DRAM[15570] = 8'b10100111;
DRAM[15571] = 8'b10101000;
DRAM[15572] = 8'b10110000;
DRAM[15573] = 8'b10111001;
DRAM[15574] = 8'b10111101;
DRAM[15575] = 8'b11000100;
DRAM[15576] = 8'b11001100;
DRAM[15577] = 8'b11010000;
DRAM[15578] = 8'b11010010;
DRAM[15579] = 8'b11010100;
DRAM[15580] = 8'b11010110;
DRAM[15581] = 8'b11010111;
DRAM[15582] = 8'b01001110;
DRAM[15583] = 8'b01100001;
DRAM[15584] = 8'b01100101;
DRAM[15585] = 8'b01100110;
DRAM[15586] = 8'b01100110;
DRAM[15587] = 8'b01100001;
DRAM[15588] = 8'b01100001;
DRAM[15589] = 8'b01010101;
DRAM[15590] = 8'b01010100;
DRAM[15591] = 8'b01010101;
DRAM[15592] = 8'b01100111;
DRAM[15593] = 8'b10110010;
DRAM[15594] = 8'b11010001;
DRAM[15595] = 8'b10111100;
DRAM[15596] = 8'b01111111;
DRAM[15597] = 8'b01001100;
DRAM[15598] = 8'b00111010;
DRAM[15599] = 8'b00111111;
DRAM[15600] = 8'b01001010;
DRAM[15601] = 8'b01000111;
DRAM[15602] = 8'b01010001;
DRAM[15603] = 8'b01100101;
DRAM[15604] = 8'b01100101;
DRAM[15605] = 8'b01011000;
DRAM[15606] = 8'b01000110;
DRAM[15607] = 8'b01001100;
DRAM[15608] = 8'b01011010;
DRAM[15609] = 8'b01101110;
DRAM[15610] = 8'b01101010;
DRAM[15611] = 8'b01011111;
DRAM[15612] = 8'b01010100;
DRAM[15613] = 8'b01000010;
DRAM[15614] = 8'b01000100;
DRAM[15615] = 8'b01000000;
DRAM[15616] = 8'b00111100;
DRAM[15617] = 8'b01011100;
DRAM[15618] = 8'b01100000;
DRAM[15619] = 8'b10000000;
DRAM[15620] = 8'b10101000;
DRAM[15621] = 8'b10110001;
DRAM[15622] = 8'b10011000;
DRAM[15623] = 8'b01011111;
DRAM[15624] = 8'b01110011;
DRAM[15625] = 8'b10011000;
DRAM[15626] = 8'b10101101;
DRAM[15627] = 8'b10110010;
DRAM[15628] = 8'b10110110;
DRAM[15629] = 8'b10110110;
DRAM[15630] = 8'b10101011;
DRAM[15631] = 8'b01111001;
DRAM[15632] = 8'b01100001;
DRAM[15633] = 8'b00101011;
DRAM[15634] = 8'b00110001;
DRAM[15635] = 8'b00110011;
DRAM[15636] = 8'b00110101;
DRAM[15637] = 8'b00111010;
DRAM[15638] = 8'b00110011;
DRAM[15639] = 8'b00110000;
DRAM[15640] = 8'b01000000;
DRAM[15641] = 8'b00110001;
DRAM[15642] = 8'b00111110;
DRAM[15643] = 8'b01011100;
DRAM[15644] = 8'b00101100;
DRAM[15645] = 8'b01001101;
DRAM[15646] = 8'b01101000;
DRAM[15647] = 8'b00111010;
DRAM[15648] = 8'b00101110;
DRAM[15649] = 8'b01010100;
DRAM[15650] = 8'b00101101;
DRAM[15651] = 8'b01010101;
DRAM[15652] = 8'b01000100;
DRAM[15653] = 8'b00111011;
DRAM[15654] = 8'b01101000;
DRAM[15655] = 8'b10000101;
DRAM[15656] = 8'b01000101;
DRAM[15657] = 8'b00111011;
DRAM[15658] = 8'b00100111;
DRAM[15659] = 8'b00110010;
DRAM[15660] = 8'b00101101;
DRAM[15661] = 8'b00101111;
DRAM[15662] = 8'b00101111;
DRAM[15663] = 8'b00110111;
DRAM[15664] = 8'b00111111;
DRAM[15665] = 8'b00101101;
DRAM[15666] = 8'b00111100;
DRAM[15667] = 8'b01001010;
DRAM[15668] = 8'b01100010;
DRAM[15669] = 8'b01101101;
DRAM[15670] = 8'b01111001;
DRAM[15671] = 8'b01111100;
DRAM[15672] = 8'b01111110;
DRAM[15673] = 8'b10000010;
DRAM[15674] = 8'b10000100;
DRAM[15675] = 8'b10001000;
DRAM[15676] = 8'b10001000;
DRAM[15677] = 8'b10001000;
DRAM[15678] = 8'b10001011;
DRAM[15679] = 8'b10001011;
DRAM[15680] = 8'b10001010;
DRAM[15681] = 8'b10001110;
DRAM[15682] = 8'b10001111;
DRAM[15683] = 8'b10001111;
DRAM[15684] = 8'b10010010;
DRAM[15685] = 8'b10010001;
DRAM[15686] = 8'b10010010;
DRAM[15687] = 8'b10001101;
DRAM[15688] = 8'b10001111;
DRAM[15689] = 8'b10001010;
DRAM[15690] = 8'b10001011;
DRAM[15691] = 8'b10001110;
DRAM[15692] = 8'b10001101;
DRAM[15693] = 8'b10010000;
DRAM[15694] = 8'b10010010;
DRAM[15695] = 8'b10010111;
DRAM[15696] = 8'b10011100;
DRAM[15697] = 8'b10011110;
DRAM[15698] = 8'b10100100;
DRAM[15699] = 8'b10101011;
DRAM[15700] = 8'b10101110;
DRAM[15701] = 8'b10110101;
DRAM[15702] = 8'b10111100;
DRAM[15703] = 8'b11000010;
DRAM[15704] = 8'b11001001;
DRAM[15705] = 8'b11001101;
DRAM[15706] = 8'b11010010;
DRAM[15707] = 8'b11010010;
DRAM[15708] = 8'b11010110;
DRAM[15709] = 8'b11010101;
DRAM[15710] = 8'b01110101;
DRAM[15711] = 8'b01011000;
DRAM[15712] = 8'b01100011;
DRAM[15713] = 8'b01100101;
DRAM[15714] = 8'b01101000;
DRAM[15715] = 8'b01100111;
DRAM[15716] = 8'b01100100;
DRAM[15717] = 8'b01100000;
DRAM[15718] = 8'b01100101;
DRAM[15719] = 8'b01100110;
DRAM[15720] = 8'b01101000;
DRAM[15721] = 8'b10011110;
DRAM[15722] = 8'b10110011;
DRAM[15723] = 8'b01111100;
DRAM[15724] = 8'b01010001;
DRAM[15725] = 8'b01001110;
DRAM[15726] = 8'b01001010;
DRAM[15727] = 8'b01001011;
DRAM[15728] = 8'b01001001;
DRAM[15729] = 8'b01010001;
DRAM[15730] = 8'b01101000;
DRAM[15731] = 8'b01101101;
DRAM[15732] = 8'b01010110;
DRAM[15733] = 8'b01001010;
DRAM[15734] = 8'b01000000;
DRAM[15735] = 8'b01010001;
DRAM[15736] = 8'b01101000;
DRAM[15737] = 8'b01110011;
DRAM[15738] = 8'b01101010;
DRAM[15739] = 8'b01011111;
DRAM[15740] = 8'b01000101;
DRAM[15741] = 8'b01000100;
DRAM[15742] = 8'b01000100;
DRAM[15743] = 8'b00110110;
DRAM[15744] = 8'b00110001;
DRAM[15745] = 8'b01000101;
DRAM[15746] = 8'b01010110;
DRAM[15747] = 8'b01110100;
DRAM[15748] = 8'b10100010;
DRAM[15749] = 8'b10101110;
DRAM[15750] = 8'b10011001;
DRAM[15751] = 8'b01101011;
DRAM[15752] = 8'b01110010;
DRAM[15753] = 8'b10010111;
DRAM[15754] = 8'b10101011;
DRAM[15755] = 8'b10110010;
DRAM[15756] = 8'b10110101;
DRAM[15757] = 8'b10111000;
DRAM[15758] = 8'b10101100;
DRAM[15759] = 8'b10000111;
DRAM[15760] = 8'b01000111;
DRAM[15761] = 8'b00101110;
DRAM[15762] = 8'b00110010;
DRAM[15763] = 8'b00110001;
DRAM[15764] = 8'b00101110;
DRAM[15765] = 8'b00111110;
DRAM[15766] = 8'b00110110;
DRAM[15767] = 8'b00110110;
DRAM[15768] = 8'b01001110;
DRAM[15769] = 8'b00101111;
DRAM[15770] = 8'b00111000;
DRAM[15771] = 8'b01010011;
DRAM[15772] = 8'b00101111;
DRAM[15773] = 8'b01001000;
DRAM[15774] = 8'b01101101;
DRAM[15775] = 8'b01010000;
DRAM[15776] = 8'b00101111;
DRAM[15777] = 8'b01011000;
DRAM[15778] = 8'b00111100;
DRAM[15779] = 8'b00110100;
DRAM[15780] = 8'b01100011;
DRAM[15781] = 8'b01000000;
DRAM[15782] = 8'b01011110;
DRAM[15783] = 8'b01101001;
DRAM[15784] = 8'b01110001;
DRAM[15785] = 8'b01000000;
DRAM[15786] = 8'b00101101;
DRAM[15787] = 8'b00110011;
DRAM[15788] = 8'b00101101;
DRAM[15789] = 8'b00101100;
DRAM[15790] = 8'b00101101;
DRAM[15791] = 8'b00110110;
DRAM[15792] = 8'b01000011;
DRAM[15793] = 8'b01010011;
DRAM[15794] = 8'b01011110;
DRAM[15795] = 8'b01101011;
DRAM[15796] = 8'b01110111;
DRAM[15797] = 8'b01111000;
DRAM[15798] = 8'b01111101;
DRAM[15799] = 8'b10000010;
DRAM[15800] = 8'b10000000;
DRAM[15801] = 8'b10000001;
DRAM[15802] = 8'b10000001;
DRAM[15803] = 8'b10000111;
DRAM[15804] = 8'b10000110;
DRAM[15805] = 8'b10001100;
DRAM[15806] = 8'b10001000;
DRAM[15807] = 8'b10001010;
DRAM[15808] = 8'b10001110;
DRAM[15809] = 8'b10001100;
DRAM[15810] = 8'b10001101;
DRAM[15811] = 8'b10010001;
DRAM[15812] = 8'b10010001;
DRAM[15813] = 8'b10010011;
DRAM[15814] = 8'b10010000;
DRAM[15815] = 8'b10010000;
DRAM[15816] = 8'b10010000;
DRAM[15817] = 8'b10001100;
DRAM[15818] = 8'b10001110;
DRAM[15819] = 8'b10001110;
DRAM[15820] = 8'b10001110;
DRAM[15821] = 8'b10001111;
DRAM[15822] = 8'b10010011;
DRAM[15823] = 8'b10010110;
DRAM[15824] = 8'b10011011;
DRAM[15825] = 8'b10011110;
DRAM[15826] = 8'b10100010;
DRAM[15827] = 8'b10100110;
DRAM[15828] = 8'b10110000;
DRAM[15829] = 8'b10110100;
DRAM[15830] = 8'b10111001;
DRAM[15831] = 8'b11000000;
DRAM[15832] = 8'b11000101;
DRAM[15833] = 8'b11001100;
DRAM[15834] = 8'b11010000;
DRAM[15835] = 8'b11010100;
DRAM[15836] = 8'b11010100;
DRAM[15837] = 8'b11010110;
DRAM[15838] = 8'b10001101;
DRAM[15839] = 8'b01010010;
DRAM[15840] = 8'b01011100;
DRAM[15841] = 8'b01100010;
DRAM[15842] = 8'b01101001;
DRAM[15843] = 8'b01101110;
DRAM[15844] = 8'b01101000;
DRAM[15845] = 8'b01101010;
DRAM[15846] = 8'b01110001;
DRAM[15847] = 8'b01110100;
DRAM[15848] = 8'b01101101;
DRAM[15849] = 8'b01110010;
DRAM[15850] = 8'b01110000;
DRAM[15851] = 8'b01011000;
DRAM[15852] = 8'b01010101;
DRAM[15853] = 8'b01011000;
DRAM[15854] = 8'b01011000;
DRAM[15855] = 8'b01001111;
DRAM[15856] = 8'b01001001;
DRAM[15857] = 8'b01100000;
DRAM[15858] = 8'b01101000;
DRAM[15859] = 8'b01011010;
DRAM[15860] = 8'b01001000;
DRAM[15861] = 8'b01000000;
DRAM[15862] = 8'b01000011;
DRAM[15863] = 8'b01100001;
DRAM[15864] = 8'b01110000;
DRAM[15865] = 8'b01110011;
DRAM[15866] = 8'b01101000;
DRAM[15867] = 8'b01011000;
DRAM[15868] = 8'b01000011;
DRAM[15869] = 8'b00111100;
DRAM[15870] = 8'b00111001;
DRAM[15871] = 8'b00110100;
DRAM[15872] = 8'b00111000;
DRAM[15873] = 8'b00111101;
DRAM[15874] = 8'b01001001;
DRAM[15875] = 8'b01100100;
DRAM[15876] = 8'b10100111;
DRAM[15877] = 8'b10111010;
DRAM[15878] = 8'b10101010;
DRAM[15879] = 8'b01110100;
DRAM[15880] = 8'b01110011;
DRAM[15881] = 8'b10010110;
DRAM[15882] = 8'b10101100;
DRAM[15883] = 8'b10110011;
DRAM[15884] = 8'b10110111;
DRAM[15885] = 8'b10110111;
DRAM[15886] = 8'b10101100;
DRAM[15887] = 8'b01101011;
DRAM[15888] = 8'b00111111;
DRAM[15889] = 8'b00111000;
DRAM[15890] = 8'b00110100;
DRAM[15891] = 8'b00110001;
DRAM[15892] = 8'b00101111;
DRAM[15893] = 8'b00111010;
DRAM[15894] = 8'b00110111;
DRAM[15895] = 8'b00111011;
DRAM[15896] = 8'b01000101;
DRAM[15897] = 8'b00101110;
DRAM[15898] = 8'b00110101;
DRAM[15899] = 8'b01001110;
DRAM[15900] = 8'b00101010;
DRAM[15901] = 8'b01001000;
DRAM[15902] = 8'b01011101;
DRAM[15903] = 8'b01110110;
DRAM[15904] = 8'b00101000;
DRAM[15905] = 8'b01010001;
DRAM[15906] = 8'b01100110;
DRAM[15907] = 8'b00100010;
DRAM[15908] = 8'b01001100;
DRAM[15909] = 8'b01010001;
DRAM[15910] = 8'b01001010;
DRAM[15911] = 8'b01110101;
DRAM[15912] = 8'b01010010;
DRAM[15913] = 8'b00111011;
DRAM[15914] = 8'b00101000;
DRAM[15915] = 8'b00110011;
DRAM[15916] = 8'b00101011;
DRAM[15917] = 8'b00110001;
DRAM[15918] = 8'b00111001;
DRAM[15919] = 8'b01010010;
DRAM[15920] = 8'b01100000;
DRAM[15921] = 8'b01101110;
DRAM[15922] = 8'b01110100;
DRAM[15923] = 8'b01110111;
DRAM[15924] = 8'b01111010;
DRAM[15925] = 8'b01111100;
DRAM[15926] = 8'b01111101;
DRAM[15927] = 8'b10000010;
DRAM[15928] = 8'b10000010;
DRAM[15929] = 8'b10000000;
DRAM[15930] = 8'b10000000;
DRAM[15931] = 8'b10000100;
DRAM[15932] = 8'b10001001;
DRAM[15933] = 8'b10000111;
DRAM[15934] = 8'b10000111;
DRAM[15935] = 8'b10001101;
DRAM[15936] = 8'b10001011;
DRAM[15937] = 8'b10001011;
DRAM[15938] = 8'b10001101;
DRAM[15939] = 8'b10001110;
DRAM[15940] = 8'b10010010;
DRAM[15941] = 8'b10010001;
DRAM[15942] = 8'b10010001;
DRAM[15943] = 8'b10010010;
DRAM[15944] = 8'b10010001;
DRAM[15945] = 8'b10010010;
DRAM[15946] = 8'b10010001;
DRAM[15947] = 8'b10010000;
DRAM[15948] = 8'b10001111;
DRAM[15949] = 8'b10010001;
DRAM[15950] = 8'b10010101;
DRAM[15951] = 8'b10010101;
DRAM[15952] = 8'b10011000;
DRAM[15953] = 8'b10011011;
DRAM[15954] = 8'b10100001;
DRAM[15955] = 8'b10100101;
DRAM[15956] = 8'b10101001;
DRAM[15957] = 8'b10110001;
DRAM[15958] = 8'b10110101;
DRAM[15959] = 8'b10111100;
DRAM[15960] = 8'b11000010;
DRAM[15961] = 8'b11000110;
DRAM[15962] = 8'b11001100;
DRAM[15963] = 8'b11010011;
DRAM[15964] = 8'b11010010;
DRAM[15965] = 8'b11010100;
DRAM[15966] = 8'b10111100;
DRAM[15967] = 8'b01001000;
DRAM[15968] = 8'b01010111;
DRAM[15969] = 8'b01100011;
DRAM[15970] = 8'b01101010;
DRAM[15971] = 8'b01101111;
DRAM[15972] = 8'b01110000;
DRAM[15973] = 8'b01110100;
DRAM[15974] = 8'b01110110;
DRAM[15975] = 8'b01110011;
DRAM[15976] = 8'b01110010;
DRAM[15977] = 8'b01101011;
DRAM[15978] = 8'b01100110;
DRAM[15979] = 8'b01011110;
DRAM[15980] = 8'b01101001;
DRAM[15981] = 8'b01101001;
DRAM[15982] = 8'b01011010;
DRAM[15983] = 8'b01010000;
DRAM[15984] = 8'b01010111;
DRAM[15985] = 8'b01100100;
DRAM[15986] = 8'b01010101;
DRAM[15987] = 8'b01001011;
DRAM[15988] = 8'b01001001;
DRAM[15989] = 8'b01000110;
DRAM[15990] = 8'b01010101;
DRAM[15991] = 8'b01101111;
DRAM[15992] = 8'b01110111;
DRAM[15993] = 8'b01101110;
DRAM[15994] = 8'b01100010;
DRAM[15995] = 8'b01001011;
DRAM[15996] = 8'b00111101;
DRAM[15997] = 8'b00111001;
DRAM[15998] = 8'b00110011;
DRAM[15999] = 8'b00110101;
DRAM[16000] = 8'b00110100;
DRAM[16001] = 8'b00110100;
DRAM[16002] = 8'b00111110;
DRAM[16003] = 8'b01100000;
DRAM[16004] = 8'b10111101;
DRAM[16005] = 8'b11001011;
DRAM[16006] = 8'b11000100;
DRAM[16007] = 8'b10000110;
DRAM[16008] = 8'b01111001;
DRAM[16009] = 8'b10010111;
DRAM[16010] = 8'b10101100;
DRAM[16011] = 8'b10110001;
DRAM[16012] = 8'b10110100;
DRAM[16013] = 8'b10110110;
DRAM[16014] = 8'b10101001;
DRAM[16015] = 8'b01101010;
DRAM[16016] = 8'b00111011;
DRAM[16017] = 8'b00110010;
DRAM[16018] = 8'b00110101;
DRAM[16019] = 8'b00110001;
DRAM[16020] = 8'b00110011;
DRAM[16021] = 8'b00111011;
DRAM[16022] = 8'b00111011;
DRAM[16023] = 8'b01000000;
DRAM[16024] = 8'b00110101;
DRAM[16025] = 8'b00111001;
DRAM[16026] = 8'b00110111;
DRAM[16027] = 8'b01101000;
DRAM[16028] = 8'b00101100;
DRAM[16029] = 8'b01010100;
DRAM[16030] = 8'b01100001;
DRAM[16031] = 8'b01110111;
DRAM[16032] = 8'b01001001;
DRAM[16033] = 8'b00110100;
DRAM[16034] = 8'b01011111;
DRAM[16035] = 8'b00111001;
DRAM[16036] = 8'b00111100;
DRAM[16037] = 8'b01011110;
DRAM[16038] = 8'b00111001;
DRAM[16039] = 8'b01010101;
DRAM[16040] = 8'b01011111;
DRAM[16041] = 8'b01001100;
DRAM[16042] = 8'b00100110;
DRAM[16043] = 8'b00110000;
DRAM[16044] = 8'b00110000;
DRAM[16045] = 8'b00111010;
DRAM[16046] = 8'b01010101;
DRAM[16047] = 8'b01100100;
DRAM[16048] = 8'b01101101;
DRAM[16049] = 8'b01110010;
DRAM[16050] = 8'b01110100;
DRAM[16051] = 8'b01110110;
DRAM[16052] = 8'b01111011;
DRAM[16053] = 8'b01111101;
DRAM[16054] = 8'b01111111;
DRAM[16055] = 8'b01111100;
DRAM[16056] = 8'b10000010;
DRAM[16057] = 8'b10000101;
DRAM[16058] = 8'b10000011;
DRAM[16059] = 8'b10000011;
DRAM[16060] = 8'b10000111;
DRAM[16061] = 8'b10000111;
DRAM[16062] = 8'b10001000;
DRAM[16063] = 8'b10001010;
DRAM[16064] = 8'b10001011;
DRAM[16065] = 8'b10001100;
DRAM[16066] = 8'b10001110;
DRAM[16067] = 8'b10001100;
DRAM[16068] = 8'b10010010;
DRAM[16069] = 8'b10010001;
DRAM[16070] = 8'b10010010;
DRAM[16071] = 8'b10010001;
DRAM[16072] = 8'b10010001;
DRAM[16073] = 8'b10010011;
DRAM[16074] = 8'b10010001;
DRAM[16075] = 8'b10010011;
DRAM[16076] = 8'b10010101;
DRAM[16077] = 8'b10010000;
DRAM[16078] = 8'b10010101;
DRAM[16079] = 8'b10010110;
DRAM[16080] = 8'b10011000;
DRAM[16081] = 8'b10011011;
DRAM[16082] = 8'b10100000;
DRAM[16083] = 8'b10100110;
DRAM[16084] = 8'b10101001;
DRAM[16085] = 8'b10101111;
DRAM[16086] = 8'b10110100;
DRAM[16087] = 8'b10111010;
DRAM[16088] = 8'b10111110;
DRAM[16089] = 8'b11000111;
DRAM[16090] = 8'b11001011;
DRAM[16091] = 8'b11001110;
DRAM[16092] = 8'b11010001;
DRAM[16093] = 8'b11010011;
DRAM[16094] = 8'b11010100;
DRAM[16095] = 8'b01001100;
DRAM[16096] = 8'b01010100;
DRAM[16097] = 8'b01100011;
DRAM[16098] = 8'b01101000;
DRAM[16099] = 8'b01101100;
DRAM[16100] = 8'b01110100;
DRAM[16101] = 8'b01110111;
DRAM[16102] = 8'b01111000;
DRAM[16103] = 8'b01110010;
DRAM[16104] = 8'b01110011;
DRAM[16105] = 8'b01101110;
DRAM[16106] = 8'b01101100;
DRAM[16107] = 8'b01101101;
DRAM[16108] = 8'b01110100;
DRAM[16109] = 8'b01101100;
DRAM[16110] = 8'b01011110;
DRAM[16111] = 8'b01011101;
DRAM[16112] = 8'b01100001;
DRAM[16113] = 8'b01011010;
DRAM[16114] = 8'b01001001;
DRAM[16115] = 8'b01001000;
DRAM[16116] = 8'b01001010;
DRAM[16117] = 8'b01010000;
DRAM[16118] = 8'b01101101;
DRAM[16119] = 8'b01111010;
DRAM[16120] = 8'b01110100;
DRAM[16121] = 8'b01100110;
DRAM[16122] = 8'b01010100;
DRAM[16123] = 8'b00111101;
DRAM[16124] = 8'b00110111;
DRAM[16125] = 8'b00111000;
DRAM[16126] = 8'b00110111;
DRAM[16127] = 8'b01000110;
DRAM[16128] = 8'b00110001;
DRAM[16129] = 8'b00110101;
DRAM[16130] = 8'b00111001;
DRAM[16131] = 8'b01011100;
DRAM[16132] = 8'b11000100;
DRAM[16133] = 8'b11001010;
DRAM[16134] = 8'b11000101;
DRAM[16135] = 8'b10011001;
DRAM[16136] = 8'b01110110;
DRAM[16137] = 8'b10011000;
DRAM[16138] = 8'b10101101;
DRAM[16139] = 8'b10101111;
DRAM[16140] = 8'b10110100;
DRAM[16141] = 8'b10110110;
DRAM[16142] = 8'b10100111;
DRAM[16143] = 8'b01101101;
DRAM[16144] = 8'b00110111;
DRAM[16145] = 8'b00110001;
DRAM[16146] = 8'b00101101;
DRAM[16147] = 8'b00110001;
DRAM[16148] = 8'b00111000;
DRAM[16149] = 8'b00111110;
DRAM[16150] = 8'b01000011;
DRAM[16151] = 8'b01000110;
DRAM[16152] = 8'b00110101;
DRAM[16153] = 8'b01001110;
DRAM[16154] = 8'b01010110;
DRAM[16155] = 8'b01001101;
DRAM[16156] = 8'b00101111;
DRAM[16157] = 8'b01010111;
DRAM[16158] = 8'b01011111;
DRAM[16159] = 8'b01001110;
DRAM[16160] = 8'b01110100;
DRAM[16161] = 8'b00101011;
DRAM[16162] = 8'b01100000;
DRAM[16163] = 8'b00111110;
DRAM[16164] = 8'b00111000;
DRAM[16165] = 8'b01010010;
DRAM[16166] = 8'b01000010;
DRAM[16167] = 8'b01000010;
DRAM[16168] = 8'b01011010;
DRAM[16169] = 8'b01110010;
DRAM[16170] = 8'b00111110;
DRAM[16171] = 8'b00100110;
DRAM[16172] = 8'b00111100;
DRAM[16173] = 8'b01001100;
DRAM[16174] = 8'b01011101;
DRAM[16175] = 8'b01101010;
DRAM[16176] = 8'b01110000;
DRAM[16177] = 8'b01110101;
DRAM[16178] = 8'b01110110;
DRAM[16179] = 8'b01111001;
DRAM[16180] = 8'b01111100;
DRAM[16181] = 8'b01111111;
DRAM[16182] = 8'b01111101;
DRAM[16183] = 8'b10000000;
DRAM[16184] = 8'b10000100;
DRAM[16185] = 8'b10000010;
DRAM[16186] = 8'b10000100;
DRAM[16187] = 8'b10000011;
DRAM[16188] = 8'b10000110;
DRAM[16189] = 8'b10001001;
DRAM[16190] = 8'b10001000;
DRAM[16191] = 8'b10001000;
DRAM[16192] = 8'b10001100;
DRAM[16193] = 8'b10001100;
DRAM[16194] = 8'b10001011;
DRAM[16195] = 8'b10001101;
DRAM[16196] = 8'b10010001;
DRAM[16197] = 8'b10010010;
DRAM[16198] = 8'b10010000;
DRAM[16199] = 8'b10010000;
DRAM[16200] = 8'b10010010;
DRAM[16201] = 8'b10010011;
DRAM[16202] = 8'b10010101;
DRAM[16203] = 8'b10010101;
DRAM[16204] = 8'b10010100;
DRAM[16205] = 8'b10010010;
DRAM[16206] = 8'b10010111;
DRAM[16207] = 8'b10011001;
DRAM[16208] = 8'b10011000;
DRAM[16209] = 8'b10011100;
DRAM[16210] = 8'b10100010;
DRAM[16211] = 8'b10100100;
DRAM[16212] = 8'b10100110;
DRAM[16213] = 8'b10101101;
DRAM[16214] = 8'b10110010;
DRAM[16215] = 8'b10111010;
DRAM[16216] = 8'b10111110;
DRAM[16217] = 8'b11000100;
DRAM[16218] = 8'b11001000;
DRAM[16219] = 8'b11001101;
DRAM[16220] = 8'b11010001;
DRAM[16221] = 8'b11010010;
DRAM[16222] = 8'b11010011;
DRAM[16223] = 8'b01110110;
DRAM[16224] = 8'b01001111;
DRAM[16225] = 8'b01011110;
DRAM[16226] = 8'b01100010;
DRAM[16227] = 8'b01101001;
DRAM[16228] = 8'b01110101;
DRAM[16229] = 8'b01110101;
DRAM[16230] = 8'b01111001;
DRAM[16231] = 8'b01111011;
DRAM[16232] = 8'b01110101;
DRAM[16233] = 8'b01110011;
DRAM[16234] = 8'b01111000;
DRAM[16235] = 8'b10000000;
DRAM[16236] = 8'b01111010;
DRAM[16237] = 8'b01100110;
DRAM[16238] = 8'b01011101;
DRAM[16239] = 8'b01100001;
DRAM[16240] = 8'b01010011;
DRAM[16241] = 8'b01010100;
DRAM[16242] = 8'b01010101;
DRAM[16243] = 8'b01001101;
DRAM[16244] = 8'b01010000;
DRAM[16245] = 8'b01101001;
DRAM[16246] = 8'b01111101;
DRAM[16247] = 8'b01111101;
DRAM[16248] = 8'b01101101;
DRAM[16249] = 8'b01011000;
DRAM[16250] = 8'b00111110;
DRAM[16251] = 8'b00110100;
DRAM[16252] = 8'b00110010;
DRAM[16253] = 8'b00111100;
DRAM[16254] = 8'b01001100;
DRAM[16255] = 8'b01011010;
DRAM[16256] = 8'b00101101;
DRAM[16257] = 8'b00110000;
DRAM[16258] = 8'b00110100;
DRAM[16259] = 8'b01010011;
DRAM[16260] = 8'b11000011;
DRAM[16261] = 8'b11000111;
DRAM[16262] = 8'b11000001;
DRAM[16263] = 8'b10010101;
DRAM[16264] = 8'b01111000;
DRAM[16265] = 8'b10010111;
DRAM[16266] = 8'b10101011;
DRAM[16267] = 8'b10110100;
DRAM[16268] = 8'b10110100;
DRAM[16269] = 8'b10110110;
DRAM[16270] = 8'b10101101;
DRAM[16271] = 8'b01010000;
DRAM[16272] = 8'b00111100;
DRAM[16273] = 8'b00101100;
DRAM[16274] = 8'b00110011;
DRAM[16275] = 8'b00110011;
DRAM[16276] = 8'b00111101;
DRAM[16277] = 8'b01000110;
DRAM[16278] = 8'b01000101;
DRAM[16279] = 8'b01000000;
DRAM[16280] = 8'b01000101;
DRAM[16281] = 8'b01001011;
DRAM[16282] = 8'b01110100;
DRAM[16283] = 8'b00110110;
DRAM[16284] = 8'b00111110;
DRAM[16285] = 8'b01011001;
DRAM[16286] = 8'b01010011;
DRAM[16287] = 8'b01010100;
DRAM[16288] = 8'b01101001;
DRAM[16289] = 8'b01001111;
DRAM[16290] = 8'b01100110;
DRAM[16291] = 8'b01000101;
DRAM[16292] = 8'b00101110;
DRAM[16293] = 8'b00111101;
DRAM[16294] = 8'b01000111;
DRAM[16295] = 8'b00110001;
DRAM[16296] = 8'b01010100;
DRAM[16297] = 8'b00111000;
DRAM[16298] = 8'b01100100;
DRAM[16299] = 8'b00111011;
DRAM[16300] = 8'b01010000;
DRAM[16301] = 8'b01010101;
DRAM[16302] = 8'b01011111;
DRAM[16303] = 8'b01101011;
DRAM[16304] = 8'b01110000;
DRAM[16305] = 8'b01110111;
DRAM[16306] = 8'b01111010;
DRAM[16307] = 8'b01111100;
DRAM[16308] = 8'b01111100;
DRAM[16309] = 8'b01111111;
DRAM[16310] = 8'b01111111;
DRAM[16311] = 8'b01111110;
DRAM[16312] = 8'b01111111;
DRAM[16313] = 8'b10000010;
DRAM[16314] = 8'b10000110;
DRAM[16315] = 8'b10000010;
DRAM[16316] = 8'b10000101;
DRAM[16317] = 8'b10001010;
DRAM[16318] = 8'b10001000;
DRAM[16319] = 8'b10000111;
DRAM[16320] = 8'b10001000;
DRAM[16321] = 8'b10001010;
DRAM[16322] = 8'b10001101;
DRAM[16323] = 8'b10001101;
DRAM[16324] = 8'b10010001;
DRAM[16325] = 8'b10010001;
DRAM[16326] = 8'b10001110;
DRAM[16327] = 8'b10010010;
DRAM[16328] = 8'b10010010;
DRAM[16329] = 8'b10010010;
DRAM[16330] = 8'b10010111;
DRAM[16331] = 8'b10010110;
DRAM[16332] = 8'b10010101;
DRAM[16333] = 8'b10010101;
DRAM[16334] = 8'b10010110;
DRAM[16335] = 8'b10010111;
DRAM[16336] = 8'b10011010;
DRAM[16337] = 8'b10011101;
DRAM[16338] = 8'b10100001;
DRAM[16339] = 8'b10100110;
DRAM[16340] = 8'b10100110;
DRAM[16341] = 8'b10101011;
DRAM[16342] = 8'b10101101;
DRAM[16343] = 8'b10110111;
DRAM[16344] = 8'b10111110;
DRAM[16345] = 8'b11000001;
DRAM[16346] = 8'b11000101;
DRAM[16347] = 8'b11001011;
DRAM[16348] = 8'b11001111;
DRAM[16349] = 8'b11010001;
DRAM[16350] = 8'b11010100;
DRAM[16351] = 8'b10011101;
DRAM[16352] = 8'b01100000;
DRAM[16353] = 8'b01011010;
DRAM[16354] = 8'b01011010;
DRAM[16355] = 8'b01100111;
DRAM[16356] = 8'b01101001;
DRAM[16357] = 8'b01111001;
DRAM[16358] = 8'b10000100;
DRAM[16359] = 8'b01111110;
DRAM[16360] = 8'b01111100;
DRAM[16361] = 8'b01111100;
DRAM[16362] = 8'b10000111;
DRAM[16363] = 8'b10000100;
DRAM[16364] = 8'b01110100;
DRAM[16365] = 8'b01011110;
DRAM[16366] = 8'b01011001;
DRAM[16367] = 8'b01001101;
DRAM[16368] = 8'b01001100;
DRAM[16369] = 8'b01011010;
DRAM[16370] = 8'b01011000;
DRAM[16371] = 8'b01010100;
DRAM[16372] = 8'b01011010;
DRAM[16373] = 8'b01110100;
DRAM[16374] = 8'b01111111;
DRAM[16375] = 8'b01111010;
DRAM[16376] = 8'b01011110;
DRAM[16377] = 8'b01000001;
DRAM[16378] = 8'b00110101;
DRAM[16379] = 8'b00101100;
DRAM[16380] = 8'b00110110;
DRAM[16381] = 8'b01000110;
DRAM[16382] = 8'b01011101;
DRAM[16383] = 8'b01100111;
end

always @ (negedge clock)
begin
    if(wren == 0)
        q <= DRAM[address];
    else
        DRAM[address] <= data;
end
endmodule